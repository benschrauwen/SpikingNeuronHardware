library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
--use IEEE.STD_LOGIC_SIGNED.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use work.utility_package.log2ceil;

entity ROM is 
	
	generic	(
	bit_lengte : integer;
	aantal_filters : integer := 88
	);
	port( 
	clk :in std_logic;
	adres_ROM : in std_logic_vector(LOG2CEIL(aantal_filters)-1 downto 0);
	A0 : out std_logic_vector(bit_lengte-1 downto 0);
	A1 : out std_logic_vector(bit_lengte-1 downto 0);
	A2 : out std_logic_vector(bit_lengte-1 downto 0);
	B0 : out std_logic_vector(bit_lengte-1 downto 0);
	B1 : out std_logic_vector(bit_lengte-1 downto 0);
	read_enable: in std_logic
	);
	
end ROM;

architecture gedrag of ROM is
type geheugen_rij is array(aantal_filters-1 downto 0) of std_logic_vector(bit_lengte-1 downto 0);

constant A0coeff :  geheugen_rij := (0=>conv_std_logic_vector(0,bit_lengte),1=>conv_std_logic_vector(13719,bit_lengte),2=>conv_std_logic_vector(14579,bit_lengte),3=>conv_std_logic_vector(14543,bit_lengte),4=>conv_std_logic_vector(14514,bit_lengte),5=>conv_std_logic_vector(14491,bit_lengte),6=>conv_std_logic_vector(14474,bit_lengte),7=>conv_std_logic_vector(14460,bit_lengte),8=>conv_std_logic_vector(14451,bit_lengte),9=>conv_std_logic_vector(14445,bit_lengte),10=>conv_std_logic_vector(14441,bit_lengte),11=>conv_std_logic_vector(14440,bit_lengte),12=>conv_std_logic_vector(14442,bit_lengte),13=>conv_std_logic_vector(14445,bit_lengte),14=>conv_std_logic_vector(14450,bit_lengte),15=>conv_std_logic_vector(14457,bit_lengte),16=>conv_std_logic_vector(14464,bit_lengte),17=>conv_std_logic_vector(14473,bit_lengte),18=>conv_std_logic_vector(14482,bit_lengte),19=>conv_std_logic_vector(14492,bit_lengte),20=>conv_std_logic_vector(14503,bit_lengte),21=>conv_std_logic_vector(14515,bit_lengte),22=>conv_std_logic_vector(14526,bit_lengte),23=>conv_std_logic_vector(14538,bit_lengte),24=>conv_std_logic_vector(14551,bit_lengte),25=>conv_std_logic_vector(14563,bit_lengte),26=>conv_std_logic_vector(14576,bit_lengte),27=>conv_std_logic_vector(14588,bit_lengte),28=>conv_std_logic_vector(14600,bit_lengte),29=>conv_std_logic_vector(14613,bit_lengte),30=>conv_std_logic_vector(14625,bit_lengte),31=>conv_std_logic_vector(14637,bit_lengte),32=>conv_std_logic_vector(14648,bit_lengte),33=>conv_std_logic_vector(14660,bit_lengte),34=>conv_std_logic_vector(14671,bit_lengte),35=>conv_std_logic_vector(14681,bit_lengte),36=>conv_std_logic_vector(14692,bit_lengte),37=>conv_std_logic_vector(14701,bit_lengte),38=>conv_std_logic_vector(14710,bit_lengte),39=>conv_std_logic_vector(14719,bit_lengte),40=>conv_std_logic_vector(14727,bit_lengte),41=>conv_std_logic_vector(14735,bit_lengte),42=>conv_std_logic_vector(14742,bit_lengte),43=>conv_std_logic_vector(14748,bit_lengte),44=>conv_std_logic_vector(14753,bit_lengte),45=>conv_std_logic_vector(14758,bit_lengte),46=>conv_std_logic_vector(14761,bit_lengte),47=>conv_std_logic_vector(14764,bit_lengte),48=>conv_std_logic_vector(14766,bit_lengte),49=>conv_std_logic_vector(14767,bit_lengte),50=>conv_std_logic_vector(14767,bit_lengte),51=>conv_std_logic_vector(14766,bit_lengte),52=>conv_std_logic_vector(14764,bit_lengte),53=>conv_std_logic_vector(14760,bit_lengte),54=>conv_std_logic_vector(14755,bit_lengte),55=>conv_std_logic_vector(14749,bit_lengte),56=>conv_std_logic_vector(14741,bit_lengte),57=>conv_std_logic_vector(14731,bit_lengte),58=>conv_std_logic_vector(14720,bit_lengte),59=>conv_std_logic_vector(14707,bit_lengte),60=>conv_std_logic_vector(14691,bit_lengte),61=>conv_std_logic_vector(14673,bit_lengte),62=>conv_std_logic_vector(14653,bit_lengte),63=>conv_std_logic_vector(14630,bit_lengte),64=>conv_std_logic_vector(14603,bit_lengte),65=>conv_std_logic_vector(14574,bit_lengte),66=>conv_std_logic_vector(14540,bit_lengte),67=>conv_std_logic_vector(14503,bit_lengte),68=>conv_std_logic_vector(14460,bit_lengte),69=>conv_std_logic_vector(14413,bit_lengte),70=>conv_std_logic_vector(14359,bit_lengte),71=>conv_std_logic_vector(14298,bit_lengte),72=>conv_std_logic_vector(14229,bit_lengte),73=>conv_std_logic_vector(14151,bit_lengte),74=>conv_std_logic_vector(14062,bit_lengte),75=>conv_std_logic_vector(13960,bit_lengte),76=>conv_std_logic_vector(13843,bit_lengte),77=>conv_std_logic_vector(13707,bit_lengte),78=>conv_std_logic_vector(13548,bit_lengte),79=>conv_std_logic_vector(13362,bit_lengte),80=>conv_std_logic_vector(13139,bit_lengte),81=>conv_std_logic_vector(12871,bit_lengte),82=>conv_std_logic_vector(12542,bit_lengte),83=>conv_std_logic_vector(12131,bit_lengte),84=>conv_std_logic_vector(11603,bit_lengte),85=>conv_std_logic_vector(10904,bit_lengte),86=>conv_std_logic_vector(9936,bit_lengte),87=>conv_std_logic_vector(8518,bit_lengte));
constant A1coeff :  geheugen_rij := (0=>conv_std_logic_vector(12246,bit_lengte),1=>conv_std_logic_vector(0,bit_lengte),2=>conv_std_logic_vector(28078,bit_lengte),3=>conv_std_logic_vector(27897,bit_lengte),4=>conv_std_logic_vector(27482,bit_lengte),5=>conv_std_logic_vector(26857,bit_lengte),6=>conv_std_logic_vector(26044,bit_lengte),7=>conv_std_logic_vector(25068,bit_lengte),8=>conv_std_logic_vector(23951,bit_lengte),9=>conv_std_logic_vector(22712,bit_lengte),10=>conv_std_logic_vector(21373,bit_lengte),11=>conv_std_logic_vector(19950,bit_lengte),12=>conv_std_logic_vector(18461,bit_lengte),13=>conv_std_logic_vector(16920,bit_lengte),14=>conv_std_logic_vector(15343,bit_lengte),15=>conv_std_logic_vector(13740,bit_lengte),16=>conv_std_logic_vector(12125,bit_lengte),17=>conv_std_logic_vector(10505,bit_lengte),18=>conv_std_logic_vector(8891,bit_lengte),19=>conv_std_logic_vector(7290,bit_lengte),20=>conv_std_logic_vector(5708,bit_lengte),21=>conv_std_logic_vector(4152,bit_lengte),22=>conv_std_logic_vector(2626,bit_lengte),23=>conv_std_logic_vector(1134,bit_lengte),24=>conv_std_logic_vector(-321,bit_lengte),25=>conv_std_logic_vector(-1736,bit_lengte),26=>conv_std_logic_vector(-3108,bit_lengte),27=>conv_std_logic_vector(-4436,bit_lengte),28=>conv_std_logic_vector(-5720,bit_lengte),29=>conv_std_logic_vector(-6958,bit_lengte),30=>conv_std_logic_vector(-8149,bit_lengte),31=>conv_std_logic_vector(-9295,bit_lengte),32=>conv_std_logic_vector(-10394,bit_lengte),33=>conv_std_logic_vector(-11448,bit_lengte),34=>conv_std_logic_vector(-12457,bit_lengte),35=>conv_std_logic_vector(-13422,bit_lengte),36=>conv_std_logic_vector(-14344,bit_lengte),37=>conv_std_logic_vector(-15223,bit_lengte),38=>conv_std_logic_vector(-16061,bit_lengte),39=>conv_std_logic_vector(-16859,bit_lengte),40=>conv_std_logic_vector(-17617,bit_lengte),41=>conv_std_logic_vector(-18339,bit_lengte),42=>conv_std_logic_vector(-19023,bit_lengte),43=>conv_std_logic_vector(-19673,bit_lengte),44=>conv_std_logic_vector(-20288,bit_lengte),45=>conv_std_logic_vector(-20870,bit_lengte),46=>conv_std_logic_vector(-21421,bit_lengte),47=>conv_std_logic_vector(-21942,bit_lengte),48=>conv_std_logic_vector(-22433,bit_lengte),49=>conv_std_logic_vector(-22897,bit_lengte),50=>conv_std_logic_vector(-23333,bit_lengte),51=>conv_std_logic_vector(-23743,bit_lengte),52=>conv_std_logic_vector(-24128,bit_lengte),53=>conv_std_logic_vector(-24489,bit_lengte),54=>conv_std_logic_vector(-24826,bit_lengte),55=>conv_std_logic_vector(-25141,bit_lengte),56=>conv_std_logic_vector(-25435,bit_lengte),57=>conv_std_logic_vector(-25707,bit_lengte),58=>conv_std_logic_vector(-25959,bit_lengte),59=>conv_std_logic_vector(-26190,bit_lengte),60=>conv_std_logic_vector(-26403,bit_lengte),61=>conv_std_logic_vector(-26596,bit_lengte),62=>conv_std_logic_vector(-26771,bit_lengte),63=>conv_std_logic_vector(-26926,bit_lengte),64=>conv_std_logic_vector(-27064,bit_lengte),65=>conv_std_logic_vector(-27183,bit_lengte),66=>conv_std_logic_vector(-27283,bit_lengte),67=>conv_std_logic_vector(-27364,bit_lengte),68=>conv_std_logic_vector(-27425,bit_lengte),69=>conv_std_logic_vector(-27466,bit_lengte),70=>conv_std_logic_vector(-27486,bit_lengte),71=>conv_std_logic_vector(-27483,bit_lengte),72=>conv_std_logic_vector(-27456,bit_lengte),73=>conv_std_logic_vector(-27402,bit_lengte),74=>conv_std_logic_vector(-27319,bit_lengte),75=>conv_std_logic_vector(-27203,bit_lengte),76=>conv_std_logic_vector(-27050,bit_lengte),77=>conv_std_logic_vector(-26853,bit_lengte),78=>conv_std_logic_vector(-26604,bit_lengte),79=>conv_std_logic_vector(-26293,bit_lengte),80=>conv_std_logic_vector(-25905,bit_lengte),81=>conv_std_logic_vector(-25420,bit_lengte),82=>conv_std_logic_vector(-24809,bit_lengte),83=>conv_std_logic_vector(-24027,bit_lengte),84=>conv_std_logic_vector(-23009,bit_lengte),85=>conv_std_logic_vector(-21643,bit_lengte),86=>conv_std_logic_vector(-19740,bit_lengte),87=>conv_std_logic_vector(-16934,bit_lengte));
constant A2coeff :  geheugen_rij := (0=>conv_std_logic_vector(-10885,bit_lengte),1=>conv_std_logic_vector(-13719,bit_lengte),2=>conv_std_logic_vector(13519,bit_lengte),3=>conv_std_logic_vector(13516,bit_lengte),4=>conv_std_logic_vector(13520,bit_lengte),5=>conv_std_logic_vector(13527,bit_lengte),6=>conv_std_logic_vector(13539,bit_lengte),7=>conv_std_logic_vector(13554,bit_lengte),8=>conv_std_logic_vector(13572,bit_lengte),9=>conv_std_logic_vector(13592,bit_lengte),10=>conv_std_logic_vector(13614,bit_lengte),11=>conv_std_logic_vector(13638,bit_lengte),12=>conv_std_logic_vector(13663,bit_lengte),13=>conv_std_logic_vector(13689,bit_lengte),14=>conv_std_logic_vector(13716,bit_lengte),15=>conv_std_logic_vector(13743,bit_lengte),16=>conv_std_logic_vector(13772,bit_lengte),17=>conv_std_logic_vector(13800,bit_lengte),18=>conv_std_logic_vector(13829,bit_lengte),19=>conv_std_logic_vector(13858,bit_lengte),20=>conv_std_logic_vector(13887,bit_lengte),21=>conv_std_logic_vector(13916,bit_lengte),22=>conv_std_logic_vector(13945,bit_lengte),23=>conv_std_logic_vector(13973,bit_lengte),24=>conv_std_logic_vector(14002,bit_lengte),25=>conv_std_logic_vector(14030,bit_lengte),26=>conv_std_logic_vector(14057,bit_lengte),27=>conv_std_logic_vector(14084,bit_lengte),28=>conv_std_logic_vector(14111,bit_lengte),29=>conv_std_logic_vector(14137,bit_lengte),30=>conv_std_logic_vector(14163,bit_lengte),31=>conv_std_logic_vector(14187,bit_lengte),32=>conv_std_logic_vector(14212,bit_lengte),33=>conv_std_logic_vector(14235,bit_lengte),34=>conv_std_logic_vector(14258,bit_lengte),35=>conv_std_logic_vector(14280,bit_lengte),36=>conv_std_logic_vector(14301,bit_lengte),37=>conv_std_logic_vector(14322,bit_lengte),38=>conv_std_logic_vector(14341,bit_lengte),39=>conv_std_logic_vector(14360,bit_lengte),40=>conv_std_logic_vector(14378,bit_lengte),41=>conv_std_logic_vector(14395,bit_lengte),42=>conv_std_logic_vector(14411,bit_lengte),43=>conv_std_logic_vector(14426,bit_lengte),44=>conv_std_logic_vector(14440,bit_lengte),45=>conv_std_logic_vector(14453,bit_lengte),46=>conv_std_logic_vector(14465,bit_lengte),47=>conv_std_logic_vector(14476,bit_lengte),48=>conv_std_logic_vector(14485,bit_lengte),49=>conv_std_logic_vector(14494,bit_lengte),50=>conv_std_logic_vector(14501,bit_lengte),51=>conv_std_logic_vector(14506,bit_lengte),52=>conv_std_logic_vector(14511,bit_lengte),53=>conv_std_logic_vector(14514,bit_lengte),54=>conv_std_logic_vector(14515,bit_lengte),55=>conv_std_logic_vector(14514,bit_lengte),56=>conv_std_logic_vector(14512,bit_lengte),57=>conv_std_logic_vector(14508,bit_lengte),58=>conv_std_logic_vector(14502,bit_lengte),59=>conv_std_logic_vector(14494,bit_lengte),60=>conv_std_logic_vector(14483,bit_lengte),61=>conv_std_logic_vector(14470,bit_lengte),62=>conv_std_logic_vector(14455,bit_lengte),63=>conv_std_logic_vector(14436,bit_lengte),64=>conv_std_logic_vector(14414,bit_lengte),65=>conv_std_logic_vector(14388,bit_lengte),66=>conv_std_logic_vector(14359,bit_lengte),67=>conv_std_logic_vector(14325,bit_lengte),68=>conv_std_logic_vector(14287,bit_lengte),69=>conv_std_logic_vector(14243,bit_lengte),70=>conv_std_logic_vector(14192,bit_lengte),71=>conv_std_logic_vector(14135,bit_lengte),72=>conv_std_logic_vector(14069,bit_lengte),73=>conv_std_logic_vector(13994,bit_lengte),74=>conv_std_logic_vector(13908,bit_lengte),75=>conv_std_logic_vector(13810,bit_lengte),76=>conv_std_logic_vector(13696,bit_lengte),77=>conv_std_logic_vector(13563,bit_lengte),78=>conv_std_logic_vector(13408,bit_lengte),79=>conv_std_logic_vector(13224,bit_lengte),80=>conv_std_logic_vector(13006,bit_lengte),81=>conv_std_logic_vector(12741,bit_lengte),82=>conv_std_logic_vector(12417,bit_lengte),83=>conv_std_logic_vector(12010,bit_lengte),84=>conv_std_logic_vector(11488,bit_lengte),85=>conv_std_logic_vector(10796,bit_lengte),86=>conv_std_logic_vector(9839,bit_lengte),87=>conv_std_logic_vector(8435,bit_lengte));
constant B0coeff :  geheugen_rij := (0=>conv_std_logic_vector(0,bit_lengte),1=>conv_std_logic_vector(26923,bit_lengte),2=>conv_std_logic_vector(26818,bit_lengte),3=>conv_std_logic_vector(26476,bit_lengte),4=>conv_std_logic_vector(25921,bit_lengte),5=>conv_std_logic_vector(25174,bit_lengte),6=>conv_std_logic_vector(24258,bit_lengte),7=>conv_std_logic_vector(23193,bit_lengte),8=>conv_std_logic_vector(21999,bit_lengte),9=>conv_std_logic_vector(20697,bit_lengte),10=>conv_std_logic_vector(19304,bit_lengte),11=>conv_std_logic_vector(17837,bit_lengte),12=>conv_std_logic_vector(16311,bit_lengte),13=>conv_std_logic_vector(14741,bit_lengte),14=>conv_std_logic_vector(13140,bit_lengte),15=>conv_std_logic_vector(11520,bit_lengte),16=>conv_std_logic_vector(9890,bit_lengte),17=>conv_std_logic_vector(8261,bit_lengte),18=>conv_std_logic_vector(6641,bit_lengte),19=>conv_std_logic_vector(5036,bit_lengte),20=>conv_std_logic_vector(3453,bit_lengte),21=>conv_std_logic_vector(1897,bit_lengte),22=>conv_std_logic_vector(372,bit_lengte),23=>conv_std_logic_vector(-1116,bit_lengte),24=>conv_std_logic_vector(-2567,bit_lengte),25=>conv_std_logic_vector(-3977,bit_lengte),26=>conv_std_logic_vector(-5344,bit_lengte),27=>conv_std_logic_vector(-6667,bit_lengte),28=>conv_std_logic_vector(-7945,bit_lengte),29=>conv_std_logic_vector(-9177,bit_lengte),30=>conv_std_logic_vector(-10364,bit_lengte),31=>conv_std_logic_vector(-11505,bit_lengte),32=>conv_std_logic_vector(-12600,bit_lengte),33=>conv_std_logic_vector(-13650,bit_lengte),34=>conv_std_logic_vector(-14656,bit_lengte),35=>conv_std_logic_vector(-15618,bit_lengte),36=>conv_std_logic_vector(-16538,bit_lengte),37=>conv_std_logic_vector(-17416,bit_lengte),38=>conv_std_logic_vector(-18254,bit_lengte),39=>conv_std_logic_vector(-19053,bit_lengte),40=>conv_std_logic_vector(-19814,bit_lengte),41=>conv_std_logic_vector(-20538,bit_lengte),42=>conv_std_logic_vector(-21227,bit_lengte),43=>conv_std_logic_vector(-21882,bit_lengte),44=>conv_std_logic_vector(-22504,bit_lengte),45=>conv_std_logic_vector(-23095,bit_lengte),46=>conv_std_logic_vector(-23655,bit_lengte),47=>conv_std_logic_vector(-24187,bit_lengte),48=>conv_std_logic_vector(-24691,bit_lengte),49=>conv_std_logic_vector(-25169,bit_lengte),50=>conv_std_logic_vector(-25621,bit_lengte),51=>conv_std_logic_vector(-26049,bit_lengte),52=>conv_std_logic_vector(-26454,bit_lengte),53=>conv_std_logic_vector(-26838,bit_lengte),54=>conv_std_logic_vector(-27200,bit_lengte),55=>conv_std_logic_vector(-27542,bit_lengte),56=>conv_std_logic_vector(-27866,bit_lengte),57=>conv_std_logic_vector(-28171,bit_lengte),58=>conv_std_logic_vector(-28459,bit_lengte),59=>conv_std_logic_vector(-28730,bit_lengte),60=>conv_std_logic_vector(-28986,bit_lengte),61=>conv_std_logic_vector(-29227,bit_lengte),62=>conv_std_logic_vector(-29454,bit_lengte),63=>conv_std_logic_vector(-29667,bit_lengte),64=>conv_std_logic_vector(-29868,bit_lengte),65=>conv_std_logic_vector(-30056,bit_lengte),66=>conv_std_logic_vector(-30233,bit_lengte),67=>conv_std_logic_vector(-30398,bit_lengte),68=>conv_std_logic_vector(-30553,bit_lengte),69=>conv_std_logic_vector(-30698,bit_lengte),70=>conv_std_logic_vector(-30833,bit_lengte),71=>conv_std_logic_vector(-30959,bit_lengte),72=>conv_std_logic_vector(-31077,bit_lengte),73=>conv_std_logic_vector(-31185,bit_lengte),74=>conv_std_logic_vector(-31286,bit_lengte),75=>conv_std_logic_vector(-31378,bit_lengte),76=>conv_std_logic_vector(-31464,bit_lengte),77=>conv_std_logic_vector(-31542,bit_lengte),78=>conv_std_logic_vector(-31613,bit_lengte),79=>conv_std_logic_vector(-31677,bit_lengte),80=>conv_std_logic_vector(-31735,bit_lengte),81=>conv_std_logic_vector(-31786,bit_lengte),82=>conv_std_logic_vector(-31831,bit_lengte),83=>conv_std_logic_vector(-31870,bit_lengte),84=>conv_std_logic_vector(-31903,bit_lengte),85=>conv_std_logic_vector(-31930,bit_lengte),86=>conv_std_logic_vector(-31952,bit_lengte),87=>conv_std_logic_vector(-31968,bit_lengte));
constant B1coeff :  geheugen_rij := (0=>conv_std_logic_vector(0,bit_lengte),1=>conv_std_logic_vector(11095,bit_lengte),2=>conv_std_logic_vector(11230,bit_lengte),3=>conv_std_logic_vector(11360,bit_lengte),4=>conv_std_logic_vector(11488,bit_lengte),5=>conv_std_logic_vector(11612,bit_lengte),6=>conv_std_logic_vector(11735,bit_lengte),7=>conv_std_logic_vector(11855,bit_lengte),8=>conv_std_logic_vector(11972,bit_lengte),9=>conv_std_logic_vector(12086,bit_lengte),10=>conv_std_logic_vector(12199,bit_lengte),11=>conv_std_logic_vector(12308,bit_lengte),12=>conv_std_logic_vector(12415,bit_lengte),13=>conv_std_logic_vector(12520,bit_lengte),14=>conv_std_logic_vector(12622,bit_lengte),15=>conv_std_logic_vector(12722,bit_lengte),16=>conv_std_logic_vector(12820,bit_lengte),17=>conv_std_logic_vector(12915,bit_lengte),18=>conv_std_logic_vector(13008,bit_lengte),19=>conv_std_logic_vector(13098,bit_lengte),20=>conv_std_logic_vector(13186,bit_lengte),21=>conv_std_logic_vector(13272,bit_lengte),22=>conv_std_logic_vector(13356,bit_lengte),23=>conv_std_logic_vector(13438,bit_lengte),24=>conv_std_logic_vector(13518,bit_lengte),25=>conv_std_logic_vector(13595,bit_lengte),26=>conv_std_logic_vector(13671,bit_lengte),27=>conv_std_logic_vector(13744,bit_lengte),28=>conv_std_logic_vector(13815,bit_lengte),29=>conv_std_logic_vector(13885,bit_lengte),30=>conv_std_logic_vector(13953,bit_lengte),31=>conv_std_logic_vector(14018,bit_lengte),32=>conv_std_logic_vector(14082,bit_lengte),33=>conv_std_logic_vector(14144,bit_lengte),34=>conv_std_logic_vector(14205,bit_lengte),35=>conv_std_logic_vector(14263,bit_lengte),36=>conv_std_logic_vector(14320,bit_lengte),37=>conv_std_logic_vector(14376,bit_lengte),38=>conv_std_logic_vector(14429,bit_lengte),39=>conv_std_logic_vector(14481,bit_lengte),40=>conv_std_logic_vector(14532,bit_lengte),41=>conv_std_logic_vector(14581,bit_lengte),42=>conv_std_logic_vector(14628,bit_lengte),43=>conv_std_logic_vector(14674,bit_lengte),44=>conv_std_logic_vector(14719,bit_lengte),45=>conv_std_logic_vector(14762,bit_lengte),46=>conv_std_logic_vector(14804,bit_lengte),47=>conv_std_logic_vector(14844,bit_lengte),48=>conv_std_logic_vector(14883,bit_lengte),49=>conv_std_logic_vector(14921,bit_lengte),50=>conv_std_logic_vector(14957,bit_lengte),51=>conv_std_logic_vector(14993,bit_lengte),52=>conv_std_logic_vector(15027,bit_lengte),53=>conv_std_logic_vector(15059,bit_lengte),54=>conv_std_logic_vector(15091,bit_lengte),55=>conv_std_logic_vector(15122,bit_lengte),56=>conv_std_logic_vector(15151,bit_lengte),57=>conv_std_logic_vector(15179,bit_lengte),58=>conv_std_logic_vector(15207,bit_lengte),59=>conv_std_logic_vector(15233,bit_lengte),60=>conv_std_logic_vector(15258,bit_lengte),61=>conv_std_logic_vector(15282,bit_lengte),62=>conv_std_logic_vector(15305,bit_lengte),63=>conv_std_logic_vector(15327,bit_lengte),64=>conv_std_logic_vector(15348,bit_lengte),65=>conv_std_logic_vector(15368,bit_lengte),66=>conv_std_logic_vector(15388,bit_lengte),67=>conv_std_logic_vector(15406,bit_lengte),68=>conv_std_logic_vector(15423,bit_lengte),69=>conv_std_logic_vector(15440,bit_lengte),70=>conv_std_logic_vector(15456,bit_lengte),71=>conv_std_logic_vector(15470,bit_lengte),72=>conv_std_logic_vector(15484,bit_lengte),73=>conv_std_logic_vector(15497,bit_lengte),74=>conv_std_logic_vector(15510,bit_lengte),75=>conv_std_logic_vector(15521,bit_lengte),76=>conv_std_logic_vector(15532,bit_lengte),77=>conv_std_logic_vector(15542,bit_lengte),78=>conv_std_logic_vector(15551,bit_lengte),79=>conv_std_logic_vector(15559,bit_lengte),80=>conv_std_logic_vector(15566,bit_lengte),81=>conv_std_logic_vector(15573,bit_lengte),82=>conv_std_logic_vector(15579,bit_lengte),83=>conv_std_logic_vector(15584,bit_lengte),84=>conv_std_logic_vector(15588,bit_lengte),85=>conv_std_logic_vector(15592,bit_lengte),86=>conv_std_logic_vector(15595,bit_lengte),87=>conv_std_logic_vector(15597,bit_lengte));

begin
	process(clk)	
	begin
		if rising_edge(clk) then
			if read_enable = '1' then --and conv_integer(adres_ROM) < aantal_filters then
				A0 <= A0coeff(conv_integer(adres_ROM));
				A1 <= A1coeff(conv_integer(adres_ROM));
				A2 <= A2coeff(conv_integer(adres_ROM));
				B0 <= B0coeff(conv_integer(adres_ROM));
				B1 <= B1coeff(conv_integer(adres_ROM));
			end if;
		end if;
	end process;
end gedrag;