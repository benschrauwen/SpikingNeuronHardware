library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_signed.all;
use work.neuron_config_package.all;
package mem_settings_package is
constant MEM : mem_type := (
conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH),
conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH),
conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(6, WEIGHT_WIDTH) & conv_std_logic_vector(3, WEIGHT_WIDTH) & conv_std_logic_vector(2, WEIGHT_WIDTH) & conv_std_logic_vector(-9, WEIGHT_WIDTH) & conv_std_logic_vector(-4, WEIGHT_WIDTH) & conv_std_logic_vector(-5, WEIGHT_WIDTH) & conv_std_logic_vector(-15, WEIGHT_WIDTH) & conv_std_logic_vector(-2, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(-18, WEIGHT_WIDTH) & conv_std_logic_vector(8, WEIGHT_WIDTH) & conv_std_logic_vector(7, WEIGHT_WIDTH) & conv_std_logic_vector(7, WEIGHT_WIDTH) & conv_std_logic_vector(-7, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(7, WEIGHT_WIDTH) & conv_std_logic_vector(6, WEIGHT_WIDTH) & conv_std_logic_vector(2, WEIGHT_WIDTH) & conv_std_logic_vector(5, WEIGHT_WIDTH) & conv_std_logic_vector(-8, WEIGHT_WIDTH) & conv_std_logic_vector(-5, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(-2, WEIGHT_WIDTH) & conv_std_logic_vector(9, WEIGHT_WIDTH) & conv_std_logic_vector(-3, WEIGHT_WIDTH) & conv_std_logic_vector(-20, WEIGHT_WIDTH) & conv_std_logic_vector(9, WEIGHT_WIDTH) & conv_std_logic_vector(-2, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(5, WEIGHT_WIDTH) & conv_std_logic_vector(2, WEIGHT_WIDTH) & conv_std_logic_vector(-4, WEIGHT_WIDTH) & conv_std_logic_vector(12, WEIGHT_WIDTH) & conv_std_logic_vector(-9, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(-8, WEIGHT_WIDTH) & conv_std_logic_vector(12, WEIGHT_WIDTH) & conv_std_logic_vector(6, WEIGHT_WIDTH) & conv_std_logic_vector(-11, WEIGHT_WIDTH) & conv_std_logic_vector(5, WEIGHT_WIDTH) & conv_std_logic_vector(-9, WEIGHT_WIDTH) & conv_std_logic_vector(-2, WEIGHT_WIDTH) & conv_std_logic_vector(3, WEIGHT_WIDTH) & conv_std_logic_vector(-7, WEIGHT_WIDTH) & conv_std_logic_vector(13, WEIGHT_WIDTH) & conv_std_logic_vector(-6, WEIGHT_WIDTH) & conv_std_logic_vector(-10, WEIGHT_WIDTH) & conv_std_logic_vector(-2, WEIGHT_WIDTH) & conv_std_logic_vector(-4, WEIGHT_WIDTH) & conv_std_logic_vector(2, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(-12, WEIGHT_WIDTH) & conv_std_logic_vector(5, WEIGHT_WIDTH) & conv_std_logic_vector(-6, WEIGHT_WIDTH) & conv_std_logic_vector(11, WEIGHT_WIDTH) & conv_std_logic_vector(-5, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(6, WEIGHT_WIDTH) & conv_std_logic_vector(-11, WEIGHT_WIDTH) & conv_std_logic_vector(4, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(15, WEIGHT_WIDTH) & conv_std_logic_vector(1, WEIGHT_WIDTH) & conv_std_logic_vector(-11, WEIGHT_WIDTH) & conv_std_logic_vector(-4, WEIGHT_WIDTH) & conv_std_logic_vector(-8, WEIGHT_WIDTH) & conv_std_logic_vector(-15, WEIGHT_WIDTH) & conv_std_logic_vector(-7, WEIGHT_WIDTH) & conv_std_logic_vector(-3, WEIGHT_WIDTH) & conv_std_logic_vector(-3, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(13, WEIGHT_WIDTH) & conv_std_logic_vector(-3, WEIGHT_WIDTH) & conv_std_logic_vector(-3, WEIGHT_WIDTH) & conv_std_logic_vector(-12, WEIGHT_WIDTH) & conv_std_logic_vector(-6, WEIGHT_WIDTH) & conv_std_logic_vector(4, WEIGHT_WIDTH) & conv_std_logic_vector(1, WEIGHT_WIDTH) & conv_std_logic_vector(-6, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(-8, WEIGHT_WIDTH) & conv_std_logic_vector(7, WEIGHT_WIDTH) & conv_std_logic_vector(13, WEIGHT_WIDTH) & conv_std_logic_vector(10, WEIGHT_WIDTH) & conv_std_logic_vector(5, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(3, WEIGHT_WIDTH) & conv_std_logic_vector(-20, WEIGHT_WIDTH) & conv_std_logic_vector(-2, WEIGHT_WIDTH) & conv_std_logic_vector(8, WEIGHT_WIDTH) & conv_std_logic_vector(3, WEIGHT_WIDTH) & conv_std_logic_vector(4, WEIGHT_WIDTH) & conv_std_logic_vector(-5, WEIGHT_WIDTH) & conv_std_logic_vector(-8, WEIGHT_WIDTH) & conv_std_logic_vector(11, WEIGHT_WIDTH) & conv_std_logic_vector(-5, WEIGHT_WIDTH) & conv_std_logic_vector(-4, WEIGHT_WIDTH) & conv_std_logic_vector(9, WEIGHT_WIDTH) & conv_std_logic_vector(12, WEIGHT_WIDTH) & conv_std_logic_vector(-5, WEIGHT_WIDTH) & conv_std_logic_vector(-12, WEIGHT_WIDTH) & conv_std_logic_vector(1, WEIGHT_WIDTH) & conv_std_logic_vector(5, WEIGHT_WIDTH) & conv_std_logic_vector(4, WEIGHT_WIDTH) & conv_std_logic_vector(2, WEIGHT_WIDTH) & conv_std_logic_vector(-12, WEIGHT_WIDTH) & conv_std_logic_vector(-7, WEIGHT_WIDTH) & conv_std_logic_vector(1, WEIGHT_WIDTH) & conv_std_logic_vector(20, WEIGHT_WIDTH) & conv_std_logic_vector(-10, WEIGHT_WIDTH) & conv_std_logic_vector(7, WEIGHT_WIDTH) & conv_std_logic_vector(-13, WEIGHT_WIDTH) & conv_std_logic_vector(13, WEIGHT_WIDTH) & conv_std_logic_vector(3, WEIGHT_WIDTH) & conv_std_logic_vector(11, WEIGHT_WIDTH) & conv_std_logic_vector(-2, WEIGHT_WIDTH) & conv_std_logic_vector(-3, WEIGHT_WIDTH) & conv_std_logic_vector(-2, WEIGHT_WIDTH) & conv_std_logic_vector(4, WEIGHT_WIDTH) & conv_std_logic_vector(-8, WEIGHT_WIDTH) & conv_std_logic_vector(18, WEIGHT_WIDTH) & conv_std_logic_vector(1, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(1, WEIGHT_WIDTH) & conv_std_logic_vector(20, WEIGHT_WIDTH) & conv_std_logic_vector(-15, WEIGHT_WIDTH) & conv_std_logic_vector(-6, WEIGHT_WIDTH) & conv_std_logic_vector(11, WEIGHT_WIDTH) & conv_std_logic_vector(-10, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(-14, WEIGHT_WIDTH) & conv_std_logic_vector(3, WEIGHT_WIDTH) & conv_std_logic_vector(-7, WEIGHT_WIDTH) & conv_std_logic_vector(4, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(11, WEIGHT_WIDTH) & conv_std_logic_vector(10, WEIGHT_WIDTH) & conv_std_logic_vector(-7, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(-6, WEIGHT_WIDTH) & conv_std_logic_vector(7, WEIGHT_WIDTH) & conv_std_logic_vector(1, WEIGHT_WIDTH) & conv_std_logic_vector(1, WEIGHT_WIDTH) & conv_std_logic_vector(2, WEIGHT_WIDTH) & conv_std_logic_vector(-2, WEIGHT_WIDTH) & conv_std_logic_vector(8, WEIGHT_WIDTH) & conv_std_logic_vector(9, WEIGHT_WIDTH) & conv_std_logic_vector(3, WEIGHT_WIDTH) & conv_std_logic_vector(-9, WEIGHT_WIDTH) & conv_std_logic_vector(-15, WEIGHT_WIDTH) & conv_std_logic_vector(12, WEIGHT_WIDTH) & conv_std_logic_vector(17, WEIGHT_WIDTH) & conv_std_logic_vector(5, WEIGHT_WIDTH) & conv_std_logic_vector(12, WEIGHT_WIDTH) & conv_std_logic_vector(9, WEIGHT_WIDTH) & conv_std_logic_vector(-10, WEIGHT_WIDTH) & conv_std_logic_vector(10, WEIGHT_WIDTH) & conv_std_logic_vector(2, WEIGHT_WIDTH) & conv_std_logic_vector(10, WEIGHT_WIDTH) & conv_std_logic_vector(-5, WEIGHT_WIDTH) & conv_std_logic_vector(1, WEIGHT_WIDTH) & conv_std_logic_vector(7, WEIGHT_WIDTH) & conv_std_logic_vector(-6, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(-10, WEIGHT_WIDTH) & conv_std_logic_vector(-9, WEIGHT_WIDTH) & conv_std_logic_vector(7, WEIGHT_WIDTH) & conv_std_logic_vector(13, WEIGHT_WIDTH) & conv_std_logic_vector(-6, WEIGHT_WIDTH) & conv_std_logic_vector(-21, WEIGHT_WIDTH) & conv_std_logic_vector(5, WEIGHT_WIDTH) & conv_std_logic_vector(-4, WEIGHT_WIDTH) & conv_std_logic_vector(-5, WEIGHT_WIDTH) & conv_std_logic_vector(1, WEIGHT_WIDTH) & conv_std_logic_vector(11, WEIGHT_WIDTH) & conv_std_logic_vector(-7, WEIGHT_WIDTH) & conv_std_logic_vector(9, WEIGHT_WIDTH) & conv_std_logic_vector(-9, WEIGHT_WIDTH) & conv_std_logic_vector(1, WEIGHT_WIDTH) & conv_std_logic_vector(6, WEIGHT_WIDTH) & conv_std_logic_vector(19, WEIGHT_WIDTH) & conv_std_logic_vector(-2, WEIGHT_WIDTH) & conv_std_logic_vector(-19, WEIGHT_WIDTH) & conv_std_logic_vector(7, WEIGHT_WIDTH) & conv_std_logic_vector(-9, WEIGHT_WIDTH) & conv_std_logic_vector(8, WEIGHT_WIDTH) & conv_std_logic_vector(-10, WEIGHT_WIDTH) & conv_std_logic_vector(3, WEIGHT_WIDTH) & conv_std_logic_vector(3, WEIGHT_WIDTH) & conv_std_logic_vector(-2, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(6, WEIGHT_WIDTH) & conv_std_logic_vector(-2, WEIGHT_WIDTH) & conv_std_logic_vector(-11, WEIGHT_WIDTH),
conv_std_logic_vector(-3, WEIGHT_WIDTH) & conv_std_logic_vector(5, WEIGHT_WIDTH) & conv_std_logic_vector(-2, WEIGHT_WIDTH) & conv_std_logic_vector(-23, WEIGHT_WIDTH) & conv_std_logic_vector(1, WEIGHT_WIDTH) & conv_std_logic_vector(10, WEIGHT_WIDTH) & conv_std_logic_vector(-10, WEIGHT_WIDTH) & conv_std_logic_vector(15, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(-5, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(1, WEIGHT_WIDTH) & conv_std_logic_vector(-21, WEIGHT_WIDTH) & conv_std_logic_vector(12, WEIGHT_WIDTH) & conv_std_logic_vector(-11, WEIGHT_WIDTH) & conv_std_logic_vector(21, WEIGHT_WIDTH) & conv_std_logic_vector(-22, WEIGHT_WIDTH) & conv_std_logic_vector(-6, WEIGHT_WIDTH) & conv_std_logic_vector(2, WEIGHT_WIDTH) & conv_std_logic_vector(-9, WEIGHT_WIDTH) & conv_std_logic_vector(18, WEIGHT_WIDTH) & conv_std_logic_vector(-12, WEIGHT_WIDTH) & conv_std_logic_vector(-13, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(6, WEIGHT_WIDTH) & conv_std_logic_vector(-6, WEIGHT_WIDTH) & conv_std_logic_vector(5, WEIGHT_WIDTH) & conv_std_logic_vector(-4, WEIGHT_WIDTH) & conv_std_logic_vector(-2, WEIGHT_WIDTH) & conv_std_logic_vector(4, WEIGHT_WIDTH) & conv_std_logic_vector(1, WEIGHT_WIDTH) & conv_std_logic_vector(-3, WEIGHT_WIDTH) & conv_std_logic_vector(14, WEIGHT_WIDTH) & conv_std_logic_vector(-9, WEIGHT_WIDTH) & conv_std_logic_vector(4, WEIGHT_WIDTH) & conv_std_logic_vector(14, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(-6, WEIGHT_WIDTH) & conv_std_logic_vector(-3, WEIGHT_WIDTH) & conv_std_logic_vector(3, WEIGHT_WIDTH) & conv_std_logic_vector(4, WEIGHT_WIDTH) & conv_std_logic_vector(6, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(2, WEIGHT_WIDTH) & conv_std_logic_vector(-9, WEIGHT_WIDTH) & conv_std_logic_vector(-6, WEIGHT_WIDTH) & conv_std_logic_vector(5, WEIGHT_WIDTH) & conv_std_logic_vector(2, WEIGHT_WIDTH) & conv_std_logic_vector(15, WEIGHT_WIDTH) & conv_std_logic_vector(-18, WEIGHT_WIDTH) & conv_std_logic_vector(10, WEIGHT_WIDTH) & conv_std_logic_vector(-7, WEIGHT_WIDTH) & conv_std_logic_vector(-5, WEIGHT_WIDTH) & conv_std_logic_vector(-8, WEIGHT_WIDTH) & conv_std_logic_vector(-2, WEIGHT_WIDTH) & conv_std_logic_vector(-4, WEIGHT_WIDTH) & conv_std_logic_vector(-11, WEIGHT_WIDTH) & conv_std_logic_vector(-7, WEIGHT_WIDTH) & conv_std_logic_vector(-9, WEIGHT_WIDTH) & conv_std_logic_vector(10, WEIGHT_WIDTH) & conv_std_logic_vector(-5, WEIGHT_WIDTH) & conv_std_logic_vector(9, WEIGHT_WIDTH) & conv_std_logic_vector(-11, WEIGHT_WIDTH) & conv_std_logic_vector(15, WEIGHT_WIDTH) & conv_std_logic_vector(9, WEIGHT_WIDTH) & conv_std_logic_vector(-4, WEIGHT_WIDTH) & conv_std_logic_vector(11, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(14, WEIGHT_WIDTH) & conv_std_logic_vector(13, WEIGHT_WIDTH) & conv_std_logic_vector(-10, WEIGHT_WIDTH) & conv_std_logic_vector(5, WEIGHT_WIDTH) & conv_std_logic_vector(4, WEIGHT_WIDTH) & conv_std_logic_vector(3, WEIGHT_WIDTH) & conv_std_logic_vector(3, WEIGHT_WIDTH) & conv_std_logic_vector(-9, WEIGHT_WIDTH) & conv_std_logic_vector(-9, WEIGHT_WIDTH) & conv_std_logic_vector(6, WEIGHT_WIDTH) & conv_std_logic_vector(2, WEIGHT_WIDTH) & conv_std_logic_vector(12, WEIGHT_WIDTH) & conv_std_logic_vector(6, WEIGHT_WIDTH) & conv_std_logic_vector(-12, WEIGHT_WIDTH) & conv_std_logic_vector(13, WEIGHT_WIDTH) & conv_std_logic_vector(-9, WEIGHT_WIDTH) & conv_std_logic_vector(8, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(3, WEIGHT_WIDTH) & conv_std_logic_vector(14, WEIGHT_WIDTH) & conv_std_logic_vector(3, WEIGHT_WIDTH) & conv_std_logic_vector(6, WEIGHT_WIDTH) & conv_std_logic_vector(5, WEIGHT_WIDTH) & conv_std_logic_vector(-2, WEIGHT_WIDTH) & conv_std_logic_vector(10, WEIGHT_WIDTH) & conv_std_logic_vector(19, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(7, WEIGHT_WIDTH) & conv_std_logic_vector(6, WEIGHT_WIDTH) & conv_std_logic_vector(3, WEIGHT_WIDTH) & conv_std_logic_vector(-11, WEIGHT_WIDTH) & conv_std_logic_vector(-10, WEIGHT_WIDTH) & conv_std_logic_vector(5, WEIGHT_WIDTH) & conv_std_logic_vector(-4, WEIGHT_WIDTH) & conv_std_logic_vector(-4, WEIGHT_WIDTH) & conv_std_logic_vector(-14, WEIGHT_WIDTH) & conv_std_logic_vector(-8, WEIGHT_WIDTH) & conv_std_logic_vector(-17, WEIGHT_WIDTH) & conv_std_logic_vector(-6, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(12, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(6, WEIGHT_WIDTH) & conv_std_logic_vector(3, WEIGHT_WIDTH) & conv_std_logic_vector(-11, WEIGHT_WIDTH) & conv_std_logic_vector(-2, WEIGHT_WIDTH) & conv_std_logic_vector(7, WEIGHT_WIDTH) & conv_std_logic_vector(-7, WEIGHT_WIDTH) & conv_std_logic_vector(-6, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(13, WEIGHT_WIDTH) & conv_std_logic_vector(-2, WEIGHT_WIDTH) & conv_std_logic_vector(-2, WEIGHT_WIDTH) & conv_std_logic_vector(1, WEIGHT_WIDTH) & conv_std_logic_vector(-19, WEIGHT_WIDTH) & conv_std_logic_vector(6, WEIGHT_WIDTH) & conv_std_logic_vector(-2, WEIGHT_WIDTH) & conv_std_logic_vector(-6, WEIGHT_WIDTH) & conv_std_logic_vector(1, WEIGHT_WIDTH) & conv_std_logic_vector(-2, WEIGHT_WIDTH) & conv_std_logic_vector(1, WEIGHT_WIDTH) & conv_std_logic_vector(8, WEIGHT_WIDTH) & conv_std_logic_vector(-22, WEIGHT_WIDTH) & conv_std_logic_vector(-16, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(2, WEIGHT_WIDTH) & conv_std_logic_vector(-6, WEIGHT_WIDTH) & conv_std_logic_vector(5, WEIGHT_WIDTH) & conv_std_logic_vector(-22, WEIGHT_WIDTH) & conv_std_logic_vector(2, WEIGHT_WIDTH) & conv_std_logic_vector(-11, WEIGHT_WIDTH) & conv_std_logic_vector(14, WEIGHT_WIDTH) & conv_std_logic_vector(9, WEIGHT_WIDTH) & conv_std_logic_vector(13, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(17, WEIGHT_WIDTH) & conv_std_logic_vector(-7, WEIGHT_WIDTH) & conv_std_logic_vector(-6, WEIGHT_WIDTH) & conv_std_logic_vector(-13, WEIGHT_WIDTH) & conv_std_logic_vector(-4, WEIGHT_WIDTH) & conv_std_logic_vector(-8, WEIGHT_WIDTH) & conv_std_logic_vector(5, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(-2, WEIGHT_WIDTH) & conv_std_logic_vector(-10, WEIGHT_WIDTH) & conv_std_logic_vector(2, WEIGHT_WIDTH) & conv_std_logic_vector(2, WEIGHT_WIDTH) & conv_std_logic_vector(2, WEIGHT_WIDTH) & conv_std_logic_vector(14, WEIGHT_WIDTH) & conv_std_logic_vector(-4, WEIGHT_WIDTH) & conv_std_logic_vector(-3, WEIGHT_WIDTH) & conv_std_logic_vector(-10, WEIGHT_WIDTH) & conv_std_logic_vector(-2, WEIGHT_WIDTH) & conv_std_logic_vector(-5, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(4, WEIGHT_WIDTH) & conv_std_logic_vector(16, WEIGHT_WIDTH) & conv_std_logic_vector(-11, WEIGHT_WIDTH) & conv_std_logic_vector(1, WEIGHT_WIDTH) & conv_std_logic_vector(-6, WEIGHT_WIDTH) & conv_std_logic_vector(1, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(-6, WEIGHT_WIDTH) & conv_std_logic_vector(-14, WEIGHT_WIDTH) & conv_std_logic_vector(-6, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(4, WEIGHT_WIDTH) & conv_std_logic_vector(2, WEIGHT_WIDTH) & conv_std_logic_vector(-11, WEIGHT_WIDTH) & conv_std_logic_vector(-13, WEIGHT_WIDTH) & conv_std_logic_vector(2, WEIGHT_WIDTH) & conv_std_logic_vector(5, WEIGHT_WIDTH) & conv_std_logic_vector(3, WEIGHT_WIDTH) & conv_std_logic_vector(-2, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(-14, WEIGHT_WIDTH) & conv_std_logic_vector(6, WEIGHT_WIDTH) & conv_std_logic_vector(-14, WEIGHT_WIDTH) & conv_std_logic_vector(11, WEIGHT_WIDTH) & conv_std_logic_vector(-15, WEIGHT_WIDTH) & conv_std_logic_vector(-11, WEIGHT_WIDTH) & conv_std_logic_vector(-5, WEIGHT_WIDTH) & conv_std_logic_vector(2, WEIGHT_WIDTH) & conv_std_logic_vector(3, WEIGHT_WIDTH) & conv_std_logic_vector(-9, WEIGHT_WIDTH) & conv_std_logic_vector(5, WEIGHT_WIDTH) & conv_std_logic_vector(-3, WEIGHT_WIDTH) & conv_std_logic_vector(3, WEIGHT_WIDTH) & conv_std_logic_vector(-7, WEIGHT_WIDTH) & conv_std_logic_vector(-8, WEIGHT_WIDTH) & conv_std_logic_vector(9, WEIGHT_WIDTH),
conv_std_logic_vector(6, WEIGHT_WIDTH) & conv_std_logic_vector(7, WEIGHT_WIDTH) & conv_std_logic_vector(2, WEIGHT_WIDTH) & conv_std_logic_vector(-14, WEIGHT_WIDTH) & conv_std_logic_vector(18, WEIGHT_WIDTH) & conv_std_logic_vector(1, WEIGHT_WIDTH) & conv_std_logic_vector(14, WEIGHT_WIDTH) & conv_std_logic_vector(1, WEIGHT_WIDTH) & conv_std_logic_vector(-3, WEIGHT_WIDTH) & conv_std_logic_vector(-7, WEIGHT_WIDTH) & conv_std_logic_vector(-12, WEIGHT_WIDTH) & conv_std_logic_vector(-2, WEIGHT_WIDTH) & conv_std_logic_vector(7, WEIGHT_WIDTH) & conv_std_logic_vector(-4, WEIGHT_WIDTH) & conv_std_logic_vector(-4, WEIGHT_WIDTH) & conv_std_logic_vector(11, WEIGHT_WIDTH) & conv_std_logic_vector(-5, WEIGHT_WIDTH) & conv_std_logic_vector(-2, WEIGHT_WIDTH) & conv_std_logic_vector(7, WEIGHT_WIDTH) & conv_std_logic_vector(14, WEIGHT_WIDTH) & conv_std_logic_vector(4, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(4, WEIGHT_WIDTH) & conv_std_logic_vector(4, WEIGHT_WIDTH) & conv_std_logic_vector(-12, WEIGHT_WIDTH) & conv_std_logic_vector(-12, WEIGHT_WIDTH) & conv_std_logic_vector(2, WEIGHT_WIDTH) & conv_std_logic_vector(5, WEIGHT_WIDTH) & conv_std_logic_vector(-5, WEIGHT_WIDTH) & conv_std_logic_vector(17, WEIGHT_WIDTH) & conv_std_logic_vector(3, WEIGHT_WIDTH) & conv_std_logic_vector(-3, WEIGHT_WIDTH) & conv_std_logic_vector(4, WEIGHT_WIDTH) & conv_std_logic_vector(-3, WEIGHT_WIDTH) & conv_std_logic_vector(5, WEIGHT_WIDTH) & conv_std_logic_vector(5, WEIGHT_WIDTH) & conv_std_logic_vector(11, WEIGHT_WIDTH) & conv_std_logic_vector(-9, WEIGHT_WIDTH) & conv_std_logic_vector(4, WEIGHT_WIDTH) & conv_std_logic_vector(-10, WEIGHT_WIDTH) & conv_std_logic_vector(-20, WEIGHT_WIDTH) & conv_std_logic_vector(-4, WEIGHT_WIDTH) & conv_std_logic_vector(2, WEIGHT_WIDTH) & conv_std_logic_vector(-2, WEIGHT_WIDTH) & conv_std_logic_vector(3, WEIGHT_WIDTH) & conv_std_logic_vector(1, WEIGHT_WIDTH) & conv_std_logic_vector(3, WEIGHT_WIDTH) & conv_std_logic_vector(3, WEIGHT_WIDTH) & conv_std_logic_vector(-17, WEIGHT_WIDTH) & conv_std_logic_vector(10, WEIGHT_WIDTH) & conv_std_logic_vector(-3, WEIGHT_WIDTH) & conv_std_logic_vector(-5, WEIGHT_WIDTH) & conv_std_logic_vector(-13, WEIGHT_WIDTH) & conv_std_logic_vector(12, WEIGHT_WIDTH) & conv_std_logic_vector(-12, WEIGHT_WIDTH) & conv_std_logic_vector(-10, WEIGHT_WIDTH) & conv_std_logic_vector(-8, WEIGHT_WIDTH) & conv_std_logic_vector(7, WEIGHT_WIDTH) & conv_std_logic_vector(2, WEIGHT_WIDTH) & conv_std_logic_vector(3, WEIGHT_WIDTH) & conv_std_logic_vector(6, WEIGHT_WIDTH) & conv_std_logic_vector(-7, WEIGHT_WIDTH) & conv_std_logic_vector(6, WEIGHT_WIDTH) & conv_std_logic_vector(3, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(-7, WEIGHT_WIDTH) & conv_std_logic_vector(12, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(17, WEIGHT_WIDTH) & conv_std_logic_vector(11, WEIGHT_WIDTH) & conv_std_logic_vector(-12, WEIGHT_WIDTH) & conv_std_logic_vector(-14, WEIGHT_WIDTH) & conv_std_logic_vector(-22, WEIGHT_WIDTH) & conv_std_logic_vector(-3, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(-13, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(-2, WEIGHT_WIDTH) & conv_std_logic_vector(1, WEIGHT_WIDTH) & conv_std_logic_vector(-2, WEIGHT_WIDTH) & conv_std_logic_vector(5, WEIGHT_WIDTH) & conv_std_logic_vector(-9, WEIGHT_WIDTH) & conv_std_logic_vector(3, WEIGHT_WIDTH) & conv_std_logic_vector(-9, WEIGHT_WIDTH) & conv_std_logic_vector(-7, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(15, WEIGHT_WIDTH) & conv_std_logic_vector(8, WEIGHT_WIDTH) & conv_std_logic_vector(-3, WEIGHT_WIDTH) & conv_std_logic_vector(13, WEIGHT_WIDTH) & conv_std_logic_vector(-3, WEIGHT_WIDTH) & conv_std_logic_vector(3, WEIGHT_WIDTH) & conv_std_logic_vector(8, WEIGHT_WIDTH) & conv_std_logic_vector(5, WEIGHT_WIDTH) & conv_std_logic_vector(-13, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(-5, WEIGHT_WIDTH) & conv_std_logic_vector(-2, WEIGHT_WIDTH) & conv_std_logic_vector(-2, WEIGHT_WIDTH) & conv_std_logic_vector(-19, WEIGHT_WIDTH) & conv_std_logic_vector(-4, WEIGHT_WIDTH) & conv_std_logic_vector(-17, WEIGHT_WIDTH) & conv_std_logic_vector(4, WEIGHT_WIDTH) & conv_std_logic_vector(1, WEIGHT_WIDTH) & conv_std_logic_vector(-3, WEIGHT_WIDTH) & conv_std_logic_vector(1, WEIGHT_WIDTH) & conv_std_logic_vector(-8, WEIGHT_WIDTH) & conv_std_logic_vector(-10, WEIGHT_WIDTH) & conv_std_logic_vector(-18, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(2, WEIGHT_WIDTH) & conv_std_logic_vector(-3, WEIGHT_WIDTH) & conv_std_logic_vector(7, WEIGHT_WIDTH) & conv_std_logic_vector(5, WEIGHT_WIDTH) & conv_std_logic_vector(-9, WEIGHT_WIDTH) & conv_std_logic_vector(7, WEIGHT_WIDTH) & conv_std_logic_vector(-16, WEIGHT_WIDTH) & conv_std_logic_vector(-2, WEIGHT_WIDTH) & conv_std_logic_vector(2, WEIGHT_WIDTH) & conv_std_logic_vector(6, WEIGHT_WIDTH) & conv_std_logic_vector(-6, WEIGHT_WIDTH) & conv_std_logic_vector(8, WEIGHT_WIDTH) & conv_std_logic_vector(-3, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(-10, WEIGHT_WIDTH) & conv_std_logic_vector(5, WEIGHT_WIDTH) & conv_std_logic_vector(2, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(3, WEIGHT_WIDTH) & conv_std_logic_vector(10, WEIGHT_WIDTH) & conv_std_logic_vector(5, WEIGHT_WIDTH) & conv_std_logic_vector(-19, WEIGHT_WIDTH) & conv_std_logic_vector(10, WEIGHT_WIDTH) & conv_std_logic_vector(-3, WEIGHT_WIDTH) & conv_std_logic_vector(-10, WEIGHT_WIDTH) & conv_std_logic_vector(12, WEIGHT_WIDTH) & conv_std_logic_vector(-6, WEIGHT_WIDTH) & conv_std_logic_vector(-3, WEIGHT_WIDTH) & conv_std_logic_vector(11, WEIGHT_WIDTH) & conv_std_logic_vector(-3, WEIGHT_WIDTH) & conv_std_logic_vector(-9, WEIGHT_WIDTH) & conv_std_logic_vector(-5, WEIGHT_WIDTH) & conv_std_logic_vector(-5, WEIGHT_WIDTH) & conv_std_logic_vector(-13, WEIGHT_WIDTH) & conv_std_logic_vector(16, WEIGHT_WIDTH) & conv_std_logic_vector(11, WEIGHT_WIDTH) & conv_std_logic_vector(-5, WEIGHT_WIDTH) & conv_std_logic_vector(-8, WEIGHT_WIDTH) & conv_std_logic_vector(-11, WEIGHT_WIDTH) & conv_std_logic_vector(-2, WEIGHT_WIDTH) & conv_std_logic_vector(-5, WEIGHT_WIDTH) & conv_std_logic_vector(-10, WEIGHT_WIDTH) & conv_std_logic_vector(17, WEIGHT_WIDTH) & conv_std_logic_vector(-16, WEIGHT_WIDTH) & conv_std_logic_vector(9, WEIGHT_WIDTH) & conv_std_logic_vector(3, WEIGHT_WIDTH) & conv_std_logic_vector(-5, WEIGHT_WIDTH) & conv_std_logic_vector(4, WEIGHT_WIDTH) & conv_std_logic_vector(-12, WEIGHT_WIDTH) & conv_std_logic_vector(-5, WEIGHT_WIDTH) & conv_std_logic_vector(7, WEIGHT_WIDTH) & conv_std_logic_vector(4, WEIGHT_WIDTH) & conv_std_logic_vector(-7, WEIGHT_WIDTH) & conv_std_logic_vector(-5, WEIGHT_WIDTH) & conv_std_logic_vector(15, WEIGHT_WIDTH) & conv_std_logic_vector(6, WEIGHT_WIDTH) & conv_std_logic_vector(4, WEIGHT_WIDTH) & conv_std_logic_vector(10, WEIGHT_WIDTH) & conv_std_logic_vector(21, WEIGHT_WIDTH) & conv_std_logic_vector(1, WEIGHT_WIDTH) & conv_std_logic_vector(3, WEIGHT_WIDTH) & conv_std_logic_vector(1, WEIGHT_WIDTH) & conv_std_logic_vector(-11, WEIGHT_WIDTH) & conv_std_logic_vector(11, WEIGHT_WIDTH) & conv_std_logic_vector(14, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(8, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(2, WEIGHT_WIDTH) & conv_std_logic_vector(13, WEIGHT_WIDTH) & conv_std_logic_vector(-13, WEIGHT_WIDTH) & conv_std_logic_vector(-6, WEIGHT_WIDTH) & conv_std_logic_vector(-6, WEIGHT_WIDTH) & conv_std_logic_vector(-8, WEIGHT_WIDTH) & conv_std_logic_vector(-9, WEIGHT_WIDTH) & conv_std_logic_vector(7, WEIGHT_WIDTH) & conv_std_logic_vector(-16, WEIGHT_WIDTH) & conv_std_logic_vector(7, WEIGHT_WIDTH) & conv_std_logic_vector(25, WEIGHT_WIDTH) & conv_std_logic_vector(-9, WEIGHT_WIDTH) & conv_std_logic_vector(-9, WEIGHT_WIDTH) & conv_std_logic_vector(1, WEIGHT_WIDTH) & conv_std_logic_vector(2, WEIGHT_WIDTH) & conv_std_logic_vector(27, WEIGHT_WIDTH) & conv_std_logic_vector(5, WEIGHT_WIDTH) & conv_std_logic_vector(6, WEIGHT_WIDTH) & conv_std_logic_vector(7, WEIGHT_WIDTH) & conv_std_logic_vector(4, WEIGHT_WIDTH) & conv_std_logic_vector(8, WEIGHT_WIDTH),
conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(-10, WEIGHT_WIDTH) & conv_std_logic_vector(-8, WEIGHT_WIDTH) & conv_std_logic_vector(8, WEIGHT_WIDTH) & conv_std_logic_vector(5, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(-13, WEIGHT_WIDTH) & conv_std_logic_vector(7, WEIGHT_WIDTH) & conv_std_logic_vector(6, WEIGHT_WIDTH) & conv_std_logic_vector(-13, WEIGHT_WIDTH) & conv_std_logic_vector(-7, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(14, WEIGHT_WIDTH) & conv_std_logic_vector(20, WEIGHT_WIDTH) & conv_std_logic_vector(2, WEIGHT_WIDTH) & conv_std_logic_vector(7, WEIGHT_WIDTH) & conv_std_logic_vector(11, WEIGHT_WIDTH) & conv_std_logic_vector(-10, WEIGHT_WIDTH) & conv_std_logic_vector(16, WEIGHT_WIDTH) & conv_std_logic_vector(-10, WEIGHT_WIDTH) & conv_std_logic_vector(10, WEIGHT_WIDTH) & conv_std_logic_vector(10, WEIGHT_WIDTH) & conv_std_logic_vector(-15, WEIGHT_WIDTH) & conv_std_logic_vector(-18, WEIGHT_WIDTH) & conv_std_logic_vector(5, WEIGHT_WIDTH) & conv_std_logic_vector(-11, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(16, WEIGHT_WIDTH) & conv_std_logic_vector(-12, WEIGHT_WIDTH) & conv_std_logic_vector(13, WEIGHT_WIDTH) & conv_std_logic_vector(-7, WEIGHT_WIDTH) & conv_std_logic_vector(20, WEIGHT_WIDTH) & conv_std_logic_vector(-3, WEIGHT_WIDTH) & conv_std_logic_vector(-18, WEIGHT_WIDTH) & conv_std_logic_vector(6, WEIGHT_WIDTH) & conv_std_logic_vector(-5, WEIGHT_WIDTH) & conv_std_logic_vector(8, WEIGHT_WIDTH) & conv_std_logic_vector(24, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(-3, WEIGHT_WIDTH) & conv_std_logic_vector(5, WEIGHT_WIDTH) & conv_std_logic_vector(-8, WEIGHT_WIDTH) & conv_std_logic_vector(-10, WEIGHT_WIDTH) & conv_std_logic_vector(2, WEIGHT_WIDTH) & conv_std_logic_vector(9, WEIGHT_WIDTH) & conv_std_logic_vector(4, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(2, WEIGHT_WIDTH) & conv_std_logic_vector(-13, WEIGHT_WIDTH) & conv_std_logic_vector(15, WEIGHT_WIDTH) & conv_std_logic_vector(-10, WEIGHT_WIDTH) & conv_std_logic_vector(-10, WEIGHT_WIDTH) & conv_std_logic_vector(-12, WEIGHT_WIDTH) & conv_std_logic_vector(-7, WEIGHT_WIDTH) & conv_std_logic_vector(-3, WEIGHT_WIDTH) & conv_std_logic_vector(1, WEIGHT_WIDTH) & conv_std_logic_vector(7, WEIGHT_WIDTH) & conv_std_logic_vector(13, WEIGHT_WIDTH) & conv_std_logic_vector(1, WEIGHT_WIDTH) & conv_std_logic_vector(9, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(4, WEIGHT_WIDTH) & conv_std_logic_vector(-13, WEIGHT_WIDTH) & conv_std_logic_vector(-11, WEIGHT_WIDTH) & conv_std_logic_vector(-4, WEIGHT_WIDTH) & conv_std_logic_vector(-24, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(-6, WEIGHT_WIDTH) & conv_std_logic_vector(-2, WEIGHT_WIDTH) & conv_std_logic_vector(-15, WEIGHT_WIDTH) & conv_std_logic_vector(24, WEIGHT_WIDTH) & conv_std_logic_vector(8, WEIGHT_WIDTH) & conv_std_logic_vector(-20, WEIGHT_WIDTH) & conv_std_logic_vector(-4, WEIGHT_WIDTH) & conv_std_logic_vector(19, WEIGHT_WIDTH) & conv_std_logic_vector(3, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(-11, WEIGHT_WIDTH) & conv_std_logic_vector(-3, WEIGHT_WIDTH) & conv_std_logic_vector(-15, WEIGHT_WIDTH) & conv_std_logic_vector(1, WEIGHT_WIDTH) & conv_std_logic_vector(-7, WEIGHT_WIDTH) & conv_std_logic_vector(1, WEIGHT_WIDTH) & conv_std_logic_vector(-8, WEIGHT_WIDTH) & conv_std_logic_vector(1, WEIGHT_WIDTH) & conv_std_logic_vector(-3, WEIGHT_WIDTH) & conv_std_logic_vector(2, WEIGHT_WIDTH) & conv_std_logic_vector(10, WEIGHT_WIDTH) & conv_std_logic_vector(14, WEIGHT_WIDTH) & conv_std_logic_vector(1, WEIGHT_WIDTH) & conv_std_logic_vector(-3, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(19, WEIGHT_WIDTH) & conv_std_logic_vector(-5, WEIGHT_WIDTH) & conv_std_logic_vector(-12, WEIGHT_WIDTH) & conv_std_logic_vector(12, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(-8, WEIGHT_WIDTH) & conv_std_logic_vector(-3, WEIGHT_WIDTH) & conv_std_logic_vector(-7, WEIGHT_WIDTH) & conv_std_logic_vector(-5, WEIGHT_WIDTH) & conv_std_logic_vector(-2, WEIGHT_WIDTH) & conv_std_logic_vector(-4, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(3, WEIGHT_WIDTH) & conv_std_logic_vector(8, WEIGHT_WIDTH) & conv_std_logic_vector(1, WEIGHT_WIDTH) & conv_std_logic_vector(-4, WEIGHT_WIDTH) & conv_std_logic_vector(-6, WEIGHT_WIDTH) & conv_std_logic_vector(-3, WEIGHT_WIDTH) & conv_std_logic_vector(-11, WEIGHT_WIDTH) & conv_std_logic_vector(-8, WEIGHT_WIDTH) & conv_std_logic_vector(10, WEIGHT_WIDTH) & conv_std_logic_vector(2, WEIGHT_WIDTH) & conv_std_logic_vector(3, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(6, WEIGHT_WIDTH) & conv_std_logic_vector(-6, WEIGHT_WIDTH) & conv_std_logic_vector(3, WEIGHT_WIDTH) & conv_std_logic_vector(-2, WEIGHT_WIDTH) & conv_std_logic_vector(-15, WEIGHT_WIDTH) & conv_std_logic_vector(7, WEIGHT_WIDTH) & conv_std_logic_vector(1, WEIGHT_WIDTH) & conv_std_logic_vector(8, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(3, WEIGHT_WIDTH) & conv_std_logic_vector(8, WEIGHT_WIDTH) & conv_std_logic_vector(-9, WEIGHT_WIDTH) & conv_std_logic_vector(-15, WEIGHT_WIDTH) & conv_std_logic_vector(4, WEIGHT_WIDTH) & conv_std_logic_vector(7, WEIGHT_WIDTH) & conv_std_logic_vector(-5, WEIGHT_WIDTH) & conv_std_logic_vector(-8, WEIGHT_WIDTH) & conv_std_logic_vector(6, WEIGHT_WIDTH) & conv_std_logic_vector(9, WEIGHT_WIDTH) & conv_std_logic_vector(16, WEIGHT_WIDTH) & conv_std_logic_vector(2, WEIGHT_WIDTH) & conv_std_logic_vector(12, WEIGHT_WIDTH) & conv_std_logic_vector(14, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(4, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(1, WEIGHT_WIDTH) & conv_std_logic_vector(12, WEIGHT_WIDTH) & conv_std_logic_vector(-8, WEIGHT_WIDTH) & conv_std_logic_vector(-5, WEIGHT_WIDTH) & conv_std_logic_vector(12, WEIGHT_WIDTH) & conv_std_logic_vector(3, WEIGHT_WIDTH) & conv_std_logic_vector(-3, WEIGHT_WIDTH) & conv_std_logic_vector(4, WEIGHT_WIDTH) & conv_std_logic_vector(-2, WEIGHT_WIDTH) & conv_std_logic_vector(16, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(8, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(4, WEIGHT_WIDTH) & conv_std_logic_vector(-3, WEIGHT_WIDTH) & conv_std_logic_vector(5, WEIGHT_WIDTH) & conv_std_logic_vector(-7, WEIGHT_WIDTH) & conv_std_logic_vector(-3, WEIGHT_WIDTH) & conv_std_logic_vector(6, WEIGHT_WIDTH) & conv_std_logic_vector(12, WEIGHT_WIDTH) & conv_std_logic_vector(-5, WEIGHT_WIDTH) & conv_std_logic_vector(-2, WEIGHT_WIDTH) & conv_std_logic_vector(9, WEIGHT_WIDTH) & conv_std_logic_vector(-7, WEIGHT_WIDTH) & conv_std_logic_vector(-9, WEIGHT_WIDTH) & conv_std_logic_vector(-5, WEIGHT_WIDTH) & conv_std_logic_vector(-5, WEIGHT_WIDTH) & conv_std_logic_vector(2, WEIGHT_WIDTH) & conv_std_logic_vector(-9, WEIGHT_WIDTH) & conv_std_logic_vector(5, WEIGHT_WIDTH) & conv_std_logic_vector(-8, WEIGHT_WIDTH) & conv_std_logic_vector(-9, WEIGHT_WIDTH) & conv_std_logic_vector(-7, WEIGHT_WIDTH) & conv_std_logic_vector(5, WEIGHT_WIDTH) & conv_std_logic_vector(6, WEIGHT_WIDTH) & conv_std_logic_vector(14, WEIGHT_WIDTH) & conv_std_logic_vector(3, WEIGHT_WIDTH) & conv_std_logic_vector(1, WEIGHT_WIDTH) & conv_std_logic_vector(-11, WEIGHT_WIDTH) & conv_std_logic_vector(-4, WEIGHT_WIDTH) & conv_std_logic_vector(12, WEIGHT_WIDTH) & conv_std_logic_vector(-19, WEIGHT_WIDTH) & conv_std_logic_vector(2, WEIGHT_WIDTH) & conv_std_logic_vector(9, WEIGHT_WIDTH) & conv_std_logic_vector(-11, WEIGHT_WIDTH) & conv_std_logic_vector(-11, WEIGHT_WIDTH) & conv_std_logic_vector(-18, WEIGHT_WIDTH) & conv_std_logic_vector(1, WEIGHT_WIDTH) & conv_std_logic_vector(-4, WEIGHT_WIDTH) & conv_std_logic_vector(-12, WEIGHT_WIDTH) & conv_std_logic_vector(7, WEIGHT_WIDTH) & conv_std_logic_vector(6, WEIGHT_WIDTH) & conv_std_logic_vector(1, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(-2, WEIGHT_WIDTH),
conv_std_logic_vector(-4, WEIGHT_WIDTH) & conv_std_logic_vector(-12, WEIGHT_WIDTH) & conv_std_logic_vector(-11, WEIGHT_WIDTH) & conv_std_logic_vector(-2, WEIGHT_WIDTH) & conv_std_logic_vector(-9, WEIGHT_WIDTH) & conv_std_logic_vector(-3, WEIGHT_WIDTH) & conv_std_logic_vector(-2, WEIGHT_WIDTH) & conv_std_logic_vector(2, WEIGHT_WIDTH) & conv_std_logic_vector(-3, WEIGHT_WIDTH) & conv_std_logic_vector(3, WEIGHT_WIDTH) & conv_std_logic_vector(-3, WEIGHT_WIDTH) & conv_std_logic_vector(-23, WEIGHT_WIDTH) & conv_std_logic_vector(1, WEIGHT_WIDTH) & conv_std_logic_vector(-7, WEIGHT_WIDTH) & conv_std_logic_vector(-2, WEIGHT_WIDTH) & conv_std_logic_vector(-13, WEIGHT_WIDTH) & conv_std_logic_vector(3, WEIGHT_WIDTH) & conv_std_logic_vector(-3, WEIGHT_WIDTH) & conv_std_logic_vector(-14, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(5, WEIGHT_WIDTH) & conv_std_logic_vector(-14, WEIGHT_WIDTH) & conv_std_logic_vector(-8, WEIGHT_WIDTH) & conv_std_logic_vector(-6, WEIGHT_WIDTH) & conv_std_logic_vector(7, WEIGHT_WIDTH) & conv_std_logic_vector(3, WEIGHT_WIDTH) & conv_std_logic_vector(6, WEIGHT_WIDTH) & conv_std_logic_vector(-2, WEIGHT_WIDTH) & conv_std_logic_vector(9, WEIGHT_WIDTH) & conv_std_logic_vector(3, WEIGHT_WIDTH) & conv_std_logic_vector(-10, WEIGHT_WIDTH) & conv_std_logic_vector(-5, WEIGHT_WIDTH) & conv_std_logic_vector(11, WEIGHT_WIDTH) & conv_std_logic_vector(-2, WEIGHT_WIDTH) & conv_std_logic_vector(11, WEIGHT_WIDTH) & conv_std_logic_vector(3, WEIGHT_WIDTH) & conv_std_logic_vector(1, WEIGHT_WIDTH) & conv_std_logic_vector(3, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(6, WEIGHT_WIDTH) & conv_std_logic_vector(17, WEIGHT_WIDTH) & conv_std_logic_vector(5, WEIGHT_WIDTH) & conv_std_logic_vector(-7, WEIGHT_WIDTH) & conv_std_logic_vector(16, WEIGHT_WIDTH) & conv_std_logic_vector(-5, WEIGHT_WIDTH) & conv_std_logic_vector(-10, WEIGHT_WIDTH) & conv_std_logic_vector(-8, WEIGHT_WIDTH) & conv_std_logic_vector(8, WEIGHT_WIDTH) & conv_std_logic_vector(-15, WEIGHT_WIDTH) & conv_std_logic_vector(5, WEIGHT_WIDTH) & conv_std_logic_vector(-10, WEIGHT_WIDTH) & conv_std_logic_vector(-2, WEIGHT_WIDTH) & conv_std_logic_vector(-14, WEIGHT_WIDTH) & conv_std_logic_vector(-5, WEIGHT_WIDTH) & conv_std_logic_vector(6, WEIGHT_WIDTH) & conv_std_logic_vector(2, WEIGHT_WIDTH) & conv_std_logic_vector(-8, WEIGHT_WIDTH) & conv_std_logic_vector(8, WEIGHT_WIDTH) & conv_std_logic_vector(8, WEIGHT_WIDTH) & conv_std_logic_vector(-13, WEIGHT_WIDTH) & conv_std_logic_vector(6, WEIGHT_WIDTH) & conv_std_logic_vector(-3, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(16, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(-5, WEIGHT_WIDTH) & conv_std_logic_vector(15, WEIGHT_WIDTH) & conv_std_logic_vector(7, WEIGHT_WIDTH) & conv_std_logic_vector(2, WEIGHT_WIDTH) & conv_std_logic_vector(5, WEIGHT_WIDTH) & conv_std_logic_vector(-6, WEIGHT_WIDTH) & conv_std_logic_vector(-4, WEIGHT_WIDTH) & conv_std_logic_vector(-6, WEIGHT_WIDTH) & conv_std_logic_vector(3, WEIGHT_WIDTH) & conv_std_logic_vector(-10, WEIGHT_WIDTH) & conv_std_logic_vector(9, WEIGHT_WIDTH) & conv_std_logic_vector(6, WEIGHT_WIDTH) & conv_std_logic_vector(-5, WEIGHT_WIDTH) & conv_std_logic_vector(10, WEIGHT_WIDTH) & conv_std_logic_vector(-4, WEIGHT_WIDTH) & conv_std_logic_vector(-14, WEIGHT_WIDTH) & conv_std_logic_vector(-11, WEIGHT_WIDTH) & conv_std_logic_vector(19, WEIGHT_WIDTH) & conv_std_logic_vector(6, WEIGHT_WIDTH) & conv_std_logic_vector(4, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(-9, WEIGHT_WIDTH) & conv_std_logic_vector(14, WEIGHT_WIDTH) & conv_std_logic_vector(-10, WEIGHT_WIDTH) & conv_std_logic_vector(7, WEIGHT_WIDTH) & conv_std_logic_vector(-19, WEIGHT_WIDTH) & conv_std_logic_vector(-11, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(-3, WEIGHT_WIDTH) & conv_std_logic_vector(-7, WEIGHT_WIDTH) & conv_std_logic_vector(-5, WEIGHT_WIDTH) & conv_std_logic_vector(8, WEIGHT_WIDTH) & conv_std_logic_vector(1, WEIGHT_WIDTH) & conv_std_logic_vector(-8, WEIGHT_WIDTH) & conv_std_logic_vector(-5, WEIGHT_WIDTH) & conv_std_logic_vector(5, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(7, WEIGHT_WIDTH) & conv_std_logic_vector(3, WEIGHT_WIDTH) & conv_std_logic_vector(-7, WEIGHT_WIDTH) & conv_std_logic_vector(-4, WEIGHT_WIDTH) & conv_std_logic_vector(7, WEIGHT_WIDTH) & conv_std_logic_vector(5, WEIGHT_WIDTH) & conv_std_logic_vector(-5, WEIGHT_WIDTH) & conv_std_logic_vector(10, WEIGHT_WIDTH) & conv_std_logic_vector(-2, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(-9, WEIGHT_WIDTH) & conv_std_logic_vector(-12, WEIGHT_WIDTH) & conv_std_logic_vector(-6, WEIGHT_WIDTH) & conv_std_logic_vector(3, WEIGHT_WIDTH) & conv_std_logic_vector(-8, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(2, WEIGHT_WIDTH) & conv_std_logic_vector(6, WEIGHT_WIDTH) & conv_std_logic_vector(5, WEIGHT_WIDTH) & conv_std_logic_vector(-12, WEIGHT_WIDTH) & conv_std_logic_vector(8, WEIGHT_WIDTH) & conv_std_logic_vector(-4, WEIGHT_WIDTH) & conv_std_logic_vector(-7, WEIGHT_WIDTH) & conv_std_logic_vector(7, WEIGHT_WIDTH) & conv_std_logic_vector(-7, WEIGHT_WIDTH) & conv_std_logic_vector(-10, WEIGHT_WIDTH) & conv_std_logic_vector(4, WEIGHT_WIDTH) & conv_std_logic_vector(1, WEIGHT_WIDTH) & conv_std_logic_vector(-20, WEIGHT_WIDTH) & conv_std_logic_vector(5, WEIGHT_WIDTH) & conv_std_logic_vector(10, WEIGHT_WIDTH) & conv_std_logic_vector(-2, WEIGHT_WIDTH) & conv_std_logic_vector(3, WEIGHT_WIDTH) & conv_std_logic_vector(9, WEIGHT_WIDTH) & conv_std_logic_vector(4, WEIGHT_WIDTH) & conv_std_logic_vector(2, WEIGHT_WIDTH) & conv_std_logic_vector(-3, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(-5, WEIGHT_WIDTH) & conv_std_logic_vector(3, WEIGHT_WIDTH) & conv_std_logic_vector(-9, WEIGHT_WIDTH) & conv_std_logic_vector(9, WEIGHT_WIDTH) & conv_std_logic_vector(2, WEIGHT_WIDTH) & conv_std_logic_vector(-4, WEIGHT_WIDTH) & conv_std_logic_vector(-4, WEIGHT_WIDTH) & conv_std_logic_vector(-4, WEIGHT_WIDTH) & conv_std_logic_vector(-9, WEIGHT_WIDTH) & conv_std_logic_vector(10, WEIGHT_WIDTH) & conv_std_logic_vector(9, WEIGHT_WIDTH) & conv_std_logic_vector(-8, WEIGHT_WIDTH) & conv_std_logic_vector(2, WEIGHT_WIDTH) & conv_std_logic_vector(4, WEIGHT_WIDTH) & conv_std_logic_vector(-6, WEIGHT_WIDTH) & conv_std_logic_vector(6, WEIGHT_WIDTH) & conv_std_logic_vector(2, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(-5, WEIGHT_WIDTH) & conv_std_logic_vector(10, WEIGHT_WIDTH) & conv_std_logic_vector(11, WEIGHT_WIDTH) & conv_std_logic_vector(-2, WEIGHT_WIDTH) & conv_std_logic_vector(-15, WEIGHT_WIDTH) & conv_std_logic_vector(2, WEIGHT_WIDTH) & conv_std_logic_vector(7, WEIGHT_WIDTH) & conv_std_logic_vector(17, WEIGHT_WIDTH) & conv_std_logic_vector(7, WEIGHT_WIDTH) & conv_std_logic_vector(1, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(-11, WEIGHT_WIDTH) & conv_std_logic_vector(13, WEIGHT_WIDTH) & conv_std_logic_vector(11, WEIGHT_WIDTH) & conv_std_logic_vector(4, WEIGHT_WIDTH) & conv_std_logic_vector(7, WEIGHT_WIDTH) & conv_std_logic_vector(5, WEIGHT_WIDTH) & conv_std_logic_vector(-2, WEIGHT_WIDTH) & conv_std_logic_vector(8, WEIGHT_WIDTH) & conv_std_logic_vector(-2, WEIGHT_WIDTH) & conv_std_logic_vector(6, WEIGHT_WIDTH) & conv_std_logic_vector(5, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(-15, WEIGHT_WIDTH) & conv_std_logic_vector(-2, WEIGHT_WIDTH) & conv_std_logic_vector(-10, WEIGHT_WIDTH) & conv_std_logic_vector(7, WEIGHT_WIDTH) & conv_std_logic_vector(11, WEIGHT_WIDTH) & conv_std_logic_vector(2, WEIGHT_WIDTH) & conv_std_logic_vector(-7, WEIGHT_WIDTH) & conv_std_logic_vector(4, WEIGHT_WIDTH) & conv_std_logic_vector(-7, WEIGHT_WIDTH) & conv_std_logic_vector(-9, WEIGHT_WIDTH) & conv_std_logic_vector(-14, WEIGHT_WIDTH) & conv_std_logic_vector(-12, WEIGHT_WIDTH) & conv_std_logic_vector(8, WEIGHT_WIDTH) & conv_std_logic_vector(-3, WEIGHT_WIDTH) & conv_std_logic_vector(6, WEIGHT_WIDTH) & conv_std_logic_vector(-2, WEIGHT_WIDTH) & conv_std_logic_vector(11, WEIGHT_WIDTH),
conv_std_logic_vector(-11, WEIGHT_WIDTH) & conv_std_logic_vector(8, WEIGHT_WIDTH) & conv_std_logic_vector(12, WEIGHT_WIDTH) & conv_std_logic_vector(5, WEIGHT_WIDTH) & conv_std_logic_vector(-9, WEIGHT_WIDTH) & conv_std_logic_vector(4, WEIGHT_WIDTH) & conv_std_logic_vector(2, WEIGHT_WIDTH) & conv_std_logic_vector(10, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(-14, WEIGHT_WIDTH) & conv_std_logic_vector(9, WEIGHT_WIDTH) & conv_std_logic_vector(3, WEIGHT_WIDTH) & conv_std_logic_vector(-9, WEIGHT_WIDTH) & conv_std_logic_vector(-5, WEIGHT_WIDTH) & conv_std_logic_vector(-6, WEIGHT_WIDTH) & conv_std_logic_vector(1, WEIGHT_WIDTH) & conv_std_logic_vector(6, WEIGHT_WIDTH) & conv_std_logic_vector(7, WEIGHT_WIDTH) & conv_std_logic_vector(-3, WEIGHT_WIDTH) & conv_std_logic_vector(-13, WEIGHT_WIDTH) & conv_std_logic_vector(3, WEIGHT_WIDTH) & conv_std_logic_vector(-13, WEIGHT_WIDTH) & conv_std_logic_vector(10, WEIGHT_WIDTH) & conv_std_logic_vector(13, WEIGHT_WIDTH) & conv_std_logic_vector(2, WEIGHT_WIDTH) & conv_std_logic_vector(-4, WEIGHT_WIDTH) & conv_std_logic_vector(2, WEIGHT_WIDTH) & conv_std_logic_vector(6, WEIGHT_WIDTH) & conv_std_logic_vector(6, WEIGHT_WIDTH) & conv_std_logic_vector(-2, WEIGHT_WIDTH) & conv_std_logic_vector(-5, WEIGHT_WIDTH) & conv_std_logic_vector(5, WEIGHT_WIDTH) & conv_std_logic_vector(-13, WEIGHT_WIDTH) & conv_std_logic_vector(3, WEIGHT_WIDTH) & conv_std_logic_vector(-11, WEIGHT_WIDTH) & conv_std_logic_vector(-3, WEIGHT_WIDTH) & conv_std_logic_vector(-8, WEIGHT_WIDTH) & conv_std_logic_vector(-8, WEIGHT_WIDTH) & conv_std_logic_vector(-10, WEIGHT_WIDTH) & conv_std_logic_vector(18, WEIGHT_WIDTH) & conv_std_logic_vector(-19, WEIGHT_WIDTH) & conv_std_logic_vector(-13, WEIGHT_WIDTH) & conv_std_logic_vector(-24, WEIGHT_WIDTH) & conv_std_logic_vector(12, WEIGHT_WIDTH) & conv_std_logic_vector(9, WEIGHT_WIDTH) & conv_std_logic_vector(-12, WEIGHT_WIDTH) & conv_std_logic_vector(17, WEIGHT_WIDTH) & conv_std_logic_vector(3, WEIGHT_WIDTH) & conv_std_logic_vector(6, WEIGHT_WIDTH) & conv_std_logic_vector(-6, WEIGHT_WIDTH) & conv_std_logic_vector(1, WEIGHT_WIDTH) & conv_std_logic_vector(-5, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(-14, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(-12, WEIGHT_WIDTH) & conv_std_logic_vector(-3, WEIGHT_WIDTH) & conv_std_logic_vector(-11, WEIGHT_WIDTH) & conv_std_logic_vector(-3, WEIGHT_WIDTH) & conv_std_logic_vector(-2, WEIGHT_WIDTH) & conv_std_logic_vector(11, WEIGHT_WIDTH) & conv_std_logic_vector(6, WEIGHT_WIDTH) & conv_std_logic_vector(2, WEIGHT_WIDTH) & conv_std_logic_vector(-8, WEIGHT_WIDTH) & conv_std_logic_vector(7, WEIGHT_WIDTH) & conv_std_logic_vector(-9, WEIGHT_WIDTH) & conv_std_logic_vector(-16, WEIGHT_WIDTH) & conv_std_logic_vector(2, WEIGHT_WIDTH) & conv_std_logic_vector(-5, WEIGHT_WIDTH) & conv_std_logic_vector(14, WEIGHT_WIDTH) & conv_std_logic_vector(3, WEIGHT_WIDTH) & conv_std_logic_vector(8, WEIGHT_WIDTH) & conv_std_logic_vector(-7, WEIGHT_WIDTH) & conv_std_logic_vector(1, WEIGHT_WIDTH) & conv_std_logic_vector(-8, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(6, WEIGHT_WIDTH) & conv_std_logic_vector(-7, WEIGHT_WIDTH) & conv_std_logic_vector(5, WEIGHT_WIDTH) & conv_std_logic_vector(4, WEIGHT_WIDTH) & conv_std_logic_vector(-7, WEIGHT_WIDTH) & conv_std_logic_vector(6, WEIGHT_WIDTH) & conv_std_logic_vector(-21, WEIGHT_WIDTH) & conv_std_logic_vector(5, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(-9, WEIGHT_WIDTH) & conv_std_logic_vector(-15, WEIGHT_WIDTH) & conv_std_logic_vector(14, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(4, WEIGHT_WIDTH) & conv_std_logic_vector(-9, WEIGHT_WIDTH) & conv_std_logic_vector(-3, WEIGHT_WIDTH) & conv_std_logic_vector(-7, WEIGHT_WIDTH) & conv_std_logic_vector(-9, WEIGHT_WIDTH) & conv_std_logic_vector(-5, WEIGHT_WIDTH) & conv_std_logic_vector(12, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(-6, WEIGHT_WIDTH) & conv_std_logic_vector(-15, WEIGHT_WIDTH) & conv_std_logic_vector(-8, WEIGHT_WIDTH) & conv_std_logic_vector(5, WEIGHT_WIDTH) & conv_std_logic_vector(-8, WEIGHT_WIDTH) & conv_std_logic_vector(-11, WEIGHT_WIDTH) & conv_std_logic_vector(-2, WEIGHT_WIDTH) & conv_std_logic_vector(13, WEIGHT_WIDTH) & conv_std_logic_vector(24, WEIGHT_WIDTH) & conv_std_logic_vector(-2, WEIGHT_WIDTH) & conv_std_logic_vector(-6, WEIGHT_WIDTH) & conv_std_logic_vector(-7, WEIGHT_WIDTH) & conv_std_logic_vector(12, WEIGHT_WIDTH) & conv_std_logic_vector(8, WEIGHT_WIDTH) & conv_std_logic_vector(8, WEIGHT_WIDTH) & conv_std_logic_vector(-3, WEIGHT_WIDTH) & conv_std_logic_vector(-6, WEIGHT_WIDTH) & conv_std_logic_vector(3, WEIGHT_WIDTH) & conv_std_logic_vector(-5, WEIGHT_WIDTH) & conv_std_logic_vector(-3, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(3, WEIGHT_WIDTH) & conv_std_logic_vector(-6, WEIGHT_WIDTH) & conv_std_logic_vector(12, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(-4, WEIGHT_WIDTH) & conv_std_logic_vector(-6, WEIGHT_WIDTH) & conv_std_logic_vector(12, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(-5, WEIGHT_WIDTH) & conv_std_logic_vector(2, WEIGHT_WIDTH) & conv_std_logic_vector(-6, WEIGHT_WIDTH) & conv_std_logic_vector(18, WEIGHT_WIDTH) & conv_std_logic_vector(-21, WEIGHT_WIDTH) & conv_std_logic_vector(-4, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(-6, WEIGHT_WIDTH) & conv_std_logic_vector(6, WEIGHT_WIDTH) & conv_std_logic_vector(-19, WEIGHT_WIDTH) & conv_std_logic_vector(6, WEIGHT_WIDTH) & conv_std_logic_vector(-7, WEIGHT_WIDTH) & conv_std_logic_vector(-16, WEIGHT_WIDTH) & conv_std_logic_vector(-6, WEIGHT_WIDTH) & conv_std_logic_vector(-5, WEIGHT_WIDTH) & conv_std_logic_vector(2, WEIGHT_WIDTH) & conv_std_logic_vector(-17, WEIGHT_WIDTH) & conv_std_logic_vector(8, WEIGHT_WIDTH) & conv_std_logic_vector(6, WEIGHT_WIDTH) & conv_std_logic_vector(4, WEIGHT_WIDTH) & conv_std_logic_vector(-5, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(-4, WEIGHT_WIDTH) & conv_std_logic_vector(11, WEIGHT_WIDTH) & conv_std_logic_vector(6, WEIGHT_WIDTH) & conv_std_logic_vector(6, WEIGHT_WIDTH) & conv_std_logic_vector(18, WEIGHT_WIDTH) & conv_std_logic_vector(7, WEIGHT_WIDTH) & conv_std_logic_vector(-9, WEIGHT_WIDTH) & conv_std_logic_vector(-15, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(1, WEIGHT_WIDTH) & conv_std_logic_vector(6, WEIGHT_WIDTH) & conv_std_logic_vector(2, WEIGHT_WIDTH) & conv_std_logic_vector(2, WEIGHT_WIDTH) & conv_std_logic_vector(-2, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(12, WEIGHT_WIDTH) & conv_std_logic_vector(-16, WEIGHT_WIDTH) & conv_std_logic_vector(-4, WEIGHT_WIDTH) & conv_std_logic_vector(3, WEIGHT_WIDTH) & conv_std_logic_vector(15, WEIGHT_WIDTH) & conv_std_logic_vector(-15, WEIGHT_WIDTH) & conv_std_logic_vector(-6, WEIGHT_WIDTH) & conv_std_logic_vector(-7, WEIGHT_WIDTH) & conv_std_logic_vector(3, WEIGHT_WIDTH) & conv_std_logic_vector(1, WEIGHT_WIDTH) & conv_std_logic_vector(8, WEIGHT_WIDTH) & conv_std_logic_vector(3, WEIGHT_WIDTH) & conv_std_logic_vector(-14, WEIGHT_WIDTH) & conv_std_logic_vector(14, WEIGHT_WIDTH) & conv_std_logic_vector(-7, WEIGHT_WIDTH) & conv_std_logic_vector(-4, WEIGHT_WIDTH) & conv_std_logic_vector(8, WEIGHT_WIDTH) & conv_std_logic_vector(-12, WEIGHT_WIDTH) & conv_std_logic_vector(3, WEIGHT_WIDTH) & conv_std_logic_vector(-5, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(-16, WEIGHT_WIDTH) & conv_std_logic_vector(8, WEIGHT_WIDTH) & conv_std_logic_vector(11, WEIGHT_WIDTH) & conv_std_logic_vector(-6, WEIGHT_WIDTH) & conv_std_logic_vector(2, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(15, WEIGHT_WIDTH) & conv_std_logic_vector(16, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(8, WEIGHT_WIDTH) & conv_std_logic_vector(-3, WEIGHT_WIDTH) & conv_std_logic_vector(-7, WEIGHT_WIDTH) & conv_std_logic_vector(-2, WEIGHT_WIDTH) & conv_std_logic_vector(2, WEIGHT_WIDTH),
conv_std_logic_vector(-4, WEIGHT_WIDTH) & conv_std_logic_vector(6, WEIGHT_WIDTH) & conv_std_logic_vector(-5, WEIGHT_WIDTH) & conv_std_logic_vector(-5, WEIGHT_WIDTH) & conv_std_logic_vector(-3, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(5, WEIGHT_WIDTH) & conv_std_logic_vector(-18, WEIGHT_WIDTH) & conv_std_logic_vector(-3, WEIGHT_WIDTH) & conv_std_logic_vector(12, WEIGHT_WIDTH) & conv_std_logic_vector(-3, WEIGHT_WIDTH) & conv_std_logic_vector(-14, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(13, WEIGHT_WIDTH) & conv_std_logic_vector(14, WEIGHT_WIDTH) & conv_std_logic_vector(6, WEIGHT_WIDTH) & conv_std_logic_vector(3, WEIGHT_WIDTH) & conv_std_logic_vector(5, WEIGHT_WIDTH) & conv_std_logic_vector(7, WEIGHT_WIDTH) & conv_std_logic_vector(5, WEIGHT_WIDTH) & conv_std_logic_vector(-6, WEIGHT_WIDTH) & conv_std_logic_vector(1, WEIGHT_WIDTH) & conv_std_logic_vector(-5, WEIGHT_WIDTH) & conv_std_logic_vector(-18, WEIGHT_WIDTH) & conv_std_logic_vector(8, WEIGHT_WIDTH) & conv_std_logic_vector(9, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(1, WEIGHT_WIDTH) & conv_std_logic_vector(-15, WEIGHT_WIDTH) & conv_std_logic_vector(-5, WEIGHT_WIDTH) & conv_std_logic_vector(15, WEIGHT_WIDTH) & conv_std_logic_vector(3, WEIGHT_WIDTH) & conv_std_logic_vector(-7, WEIGHT_WIDTH) & conv_std_logic_vector(-17, WEIGHT_WIDTH) & conv_std_logic_vector(-4, WEIGHT_WIDTH) & conv_std_logic_vector(2, WEIGHT_WIDTH) & conv_std_logic_vector(-2, WEIGHT_WIDTH) & conv_std_logic_vector(12, WEIGHT_WIDTH) & conv_std_logic_vector(-4, WEIGHT_WIDTH) & conv_std_logic_vector(4, WEIGHT_WIDTH) & conv_std_logic_vector(-2, WEIGHT_WIDTH) & conv_std_logic_vector(9, WEIGHT_WIDTH) & conv_std_logic_vector(-7, WEIGHT_WIDTH) & conv_std_logic_vector(-19, WEIGHT_WIDTH) & conv_std_logic_vector(-15, WEIGHT_WIDTH) & conv_std_logic_vector(14, WEIGHT_WIDTH) & conv_std_logic_vector(9, WEIGHT_WIDTH) & conv_std_logic_vector(21, WEIGHT_WIDTH) & conv_std_logic_vector(19, WEIGHT_WIDTH) & conv_std_logic_vector(-27, WEIGHT_WIDTH) & conv_std_logic_vector(-2, WEIGHT_WIDTH) & conv_std_logic_vector(-13, WEIGHT_WIDTH) & conv_std_logic_vector(6, WEIGHT_WIDTH) & conv_std_logic_vector(-14, WEIGHT_WIDTH) & conv_std_logic_vector(19, WEIGHT_WIDTH) & conv_std_logic_vector(2, WEIGHT_WIDTH) & conv_std_logic_vector(-7, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(-17, WEIGHT_WIDTH) & conv_std_logic_vector(7, WEIGHT_WIDTH) & conv_std_logic_vector(-5, WEIGHT_WIDTH) & conv_std_logic_vector(-5, WEIGHT_WIDTH) & conv_std_logic_vector(3, WEIGHT_WIDTH) & conv_std_logic_vector(2, WEIGHT_WIDTH) & conv_std_logic_vector(16, WEIGHT_WIDTH) & conv_std_logic_vector(-3, WEIGHT_WIDTH) & conv_std_logic_vector(-13, WEIGHT_WIDTH) & conv_std_logic_vector(13, WEIGHT_WIDTH) & conv_std_logic_vector(6, WEIGHT_WIDTH) & conv_std_logic_vector(4, WEIGHT_WIDTH) & conv_std_logic_vector(8, WEIGHT_WIDTH) & conv_std_logic_vector(-13, WEIGHT_WIDTH) & conv_std_logic_vector(-4, WEIGHT_WIDTH) & conv_std_logic_vector(8, WEIGHT_WIDTH) & conv_std_logic_vector(29, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(2, WEIGHT_WIDTH) & conv_std_logic_vector(-23, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(1, WEIGHT_WIDTH) & conv_std_logic_vector(4, WEIGHT_WIDTH) & conv_std_logic_vector(14, WEIGHT_WIDTH) & conv_std_logic_vector(-14, WEIGHT_WIDTH) & conv_std_logic_vector(6, WEIGHT_WIDTH) & conv_std_logic_vector(4, WEIGHT_WIDTH) & conv_std_logic_vector(-9, WEIGHT_WIDTH) & conv_std_logic_vector(-5, WEIGHT_WIDTH) & conv_std_logic_vector(13, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(-15, WEIGHT_WIDTH) & conv_std_logic_vector(12, WEIGHT_WIDTH) & conv_std_logic_vector(-4, WEIGHT_WIDTH) & conv_std_logic_vector(11, WEIGHT_WIDTH) & conv_std_logic_vector(20, WEIGHT_WIDTH) & conv_std_logic_vector(-22, WEIGHT_WIDTH) & conv_std_logic_vector(7, WEIGHT_WIDTH) & conv_std_logic_vector(-18, WEIGHT_WIDTH) & conv_std_logic_vector(-20, WEIGHT_WIDTH) & conv_std_logic_vector(14, WEIGHT_WIDTH) & conv_std_logic_vector(2, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(7, WEIGHT_WIDTH) & conv_std_logic_vector(-10, WEIGHT_WIDTH) & conv_std_logic_vector(8, WEIGHT_WIDTH) & conv_std_logic_vector(10, WEIGHT_WIDTH) & conv_std_logic_vector(1, WEIGHT_WIDTH) & conv_std_logic_vector(-16, WEIGHT_WIDTH) & conv_std_logic_vector(11, WEIGHT_WIDTH) & conv_std_logic_vector(-8, WEIGHT_WIDTH) & conv_std_logic_vector(18, WEIGHT_WIDTH) & conv_std_logic_vector(-3, WEIGHT_WIDTH) & conv_std_logic_vector(-10, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(4, WEIGHT_WIDTH) & conv_std_logic_vector(7, WEIGHT_WIDTH) & conv_std_logic_vector(-6, WEIGHT_WIDTH) & conv_std_logic_vector(-12, WEIGHT_WIDTH) & conv_std_logic_vector(-10, WEIGHT_WIDTH) & conv_std_logic_vector(-7, WEIGHT_WIDTH) & conv_std_logic_vector(-21, WEIGHT_WIDTH) & conv_std_logic_vector(5, WEIGHT_WIDTH) & conv_std_logic_vector(-5, WEIGHT_WIDTH) & conv_std_logic_vector(15, WEIGHT_WIDTH) & conv_std_logic_vector(-12, WEIGHT_WIDTH) & conv_std_logic_vector(21, WEIGHT_WIDTH) & conv_std_logic_vector(-9, WEIGHT_WIDTH) & conv_std_logic_vector(12, WEIGHT_WIDTH) & conv_std_logic_vector(6, WEIGHT_WIDTH) & conv_std_logic_vector(-15, WEIGHT_WIDTH) & conv_std_logic_vector(1, WEIGHT_WIDTH) & conv_std_logic_vector(4, WEIGHT_WIDTH) & conv_std_logic_vector(7, WEIGHT_WIDTH) & conv_std_logic_vector(5, WEIGHT_WIDTH) & conv_std_logic_vector(-4, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(7, WEIGHT_WIDTH) & conv_std_logic_vector(-14, WEIGHT_WIDTH) & conv_std_logic_vector(3, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(-4, WEIGHT_WIDTH) & conv_std_logic_vector(7, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(9, WEIGHT_WIDTH) & conv_std_logic_vector(9, WEIGHT_WIDTH) & conv_std_logic_vector(4, WEIGHT_WIDTH) & conv_std_logic_vector(7, WEIGHT_WIDTH) & conv_std_logic_vector(3, WEIGHT_WIDTH) & conv_std_logic_vector(5, WEIGHT_WIDTH) & conv_std_logic_vector(-4, WEIGHT_WIDTH) & conv_std_logic_vector(10, WEIGHT_WIDTH) & conv_std_logic_vector(4, WEIGHT_WIDTH) & conv_std_logic_vector(1, WEIGHT_WIDTH) & conv_std_logic_vector(-7, WEIGHT_WIDTH) & conv_std_logic_vector(4, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(-16, WEIGHT_WIDTH) & conv_std_logic_vector(2, WEIGHT_WIDTH) & conv_std_logic_vector(-13, WEIGHT_WIDTH) & conv_std_logic_vector(5, WEIGHT_WIDTH) & conv_std_logic_vector(12, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(-12, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(9, WEIGHT_WIDTH) & conv_std_logic_vector(23, WEIGHT_WIDTH) & conv_std_logic_vector(8, WEIGHT_WIDTH) & conv_std_logic_vector(-13, WEIGHT_WIDTH) & conv_std_logic_vector(2, WEIGHT_WIDTH) & conv_std_logic_vector(10, WEIGHT_WIDTH) & conv_std_logic_vector(14, WEIGHT_WIDTH) & conv_std_logic_vector(12, WEIGHT_WIDTH) & conv_std_logic_vector(12, WEIGHT_WIDTH) & conv_std_logic_vector(6, WEIGHT_WIDTH) & conv_std_logic_vector(6, WEIGHT_WIDTH) & conv_std_logic_vector(2, WEIGHT_WIDTH) & conv_std_logic_vector(2, WEIGHT_WIDTH) & conv_std_logic_vector(-16, WEIGHT_WIDTH) & conv_std_logic_vector(2, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(-5, WEIGHT_WIDTH) & conv_std_logic_vector(3, WEIGHT_WIDTH) & conv_std_logic_vector(-8, WEIGHT_WIDTH) & conv_std_logic_vector(2, WEIGHT_WIDTH) & conv_std_logic_vector(13, WEIGHT_WIDTH) & conv_std_logic_vector(12, WEIGHT_WIDTH) & conv_std_logic_vector(7, WEIGHT_WIDTH) & conv_std_logic_vector(4, WEIGHT_WIDTH) & conv_std_logic_vector(-19, WEIGHT_WIDTH) & conv_std_logic_vector(3, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(-8, WEIGHT_WIDTH) & conv_std_logic_vector(12, WEIGHT_WIDTH) & conv_std_logic_vector(11, WEIGHT_WIDTH) & conv_std_logic_vector(1, WEIGHT_WIDTH) & conv_std_logic_vector(-13, WEIGHT_WIDTH) & conv_std_logic_vector(-5, WEIGHT_WIDTH) & conv_std_logic_vector(-12, WEIGHT_WIDTH) & conv_std_logic_vector(-13, WEIGHT_WIDTH) & conv_std_logic_vector(-7, WEIGHT_WIDTH),
conv_std_logic_vector(12, WEIGHT_WIDTH) & conv_std_logic_vector(-9, WEIGHT_WIDTH) & conv_std_logic_vector(14, WEIGHT_WIDTH) & conv_std_logic_vector(7, WEIGHT_WIDTH) & conv_std_logic_vector(1, WEIGHT_WIDTH) & conv_std_logic_vector(7, WEIGHT_WIDTH) & conv_std_logic_vector(6, WEIGHT_WIDTH) & conv_std_logic_vector(-8, WEIGHT_WIDTH) & conv_std_logic_vector(7, WEIGHT_WIDTH) & conv_std_logic_vector(3, WEIGHT_WIDTH) & conv_std_logic_vector(-2, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(18, WEIGHT_WIDTH) & conv_std_logic_vector(-4, WEIGHT_WIDTH) & conv_std_logic_vector(-2, WEIGHT_WIDTH) & conv_std_logic_vector(3, WEIGHT_WIDTH) & conv_std_logic_vector(5, WEIGHT_WIDTH) & conv_std_logic_vector(1, WEIGHT_WIDTH) & conv_std_logic_vector(12, WEIGHT_WIDTH) & conv_std_logic_vector(-5, WEIGHT_WIDTH) & conv_std_logic_vector(3, WEIGHT_WIDTH) & conv_std_logic_vector(-6, WEIGHT_WIDTH) & conv_std_logic_vector(2, WEIGHT_WIDTH) & conv_std_logic_vector(-8, WEIGHT_WIDTH) & conv_std_logic_vector(7, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(-16, WEIGHT_WIDTH) & conv_std_logic_vector(2, WEIGHT_WIDTH) & conv_std_logic_vector(-9, WEIGHT_WIDTH) & conv_std_logic_vector(6, WEIGHT_WIDTH) & conv_std_logic_vector(2, WEIGHT_WIDTH) & conv_std_logic_vector(10, WEIGHT_WIDTH) & conv_std_logic_vector(9, WEIGHT_WIDTH) & conv_std_logic_vector(2, WEIGHT_WIDTH) & conv_std_logic_vector(-17, WEIGHT_WIDTH) & conv_std_logic_vector(-4, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(17, WEIGHT_WIDTH) & conv_std_logic_vector(-15, WEIGHT_WIDTH) & conv_std_logic_vector(-5, WEIGHT_WIDTH) & conv_std_logic_vector(4, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(3, WEIGHT_WIDTH) & conv_std_logic_vector(-7, WEIGHT_WIDTH) & conv_std_logic_vector(9, WEIGHT_WIDTH) & conv_std_logic_vector(6, WEIGHT_WIDTH) & conv_std_logic_vector(13, WEIGHT_WIDTH) & conv_std_logic_vector(4, WEIGHT_WIDTH) & conv_std_logic_vector(-17, WEIGHT_WIDTH) & conv_std_logic_vector(5, WEIGHT_WIDTH) & conv_std_logic_vector(5, WEIGHT_WIDTH) & conv_std_logic_vector(2, WEIGHT_WIDTH) & conv_std_logic_vector(1, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(5, WEIGHT_WIDTH) & conv_std_logic_vector(-12, WEIGHT_WIDTH) & conv_std_logic_vector(-5, WEIGHT_WIDTH) & conv_std_logic_vector(11, WEIGHT_WIDTH) & conv_std_logic_vector(-6, WEIGHT_WIDTH) & conv_std_logic_vector(-5, WEIGHT_WIDTH) & conv_std_logic_vector(-5, WEIGHT_WIDTH) & conv_std_logic_vector(-2, WEIGHT_WIDTH) & conv_std_logic_vector(19, WEIGHT_WIDTH) & conv_std_logic_vector(2, WEIGHT_WIDTH) & conv_std_logic_vector(1, WEIGHT_WIDTH) & conv_std_logic_vector(16, WEIGHT_WIDTH) & conv_std_logic_vector(-3, WEIGHT_WIDTH) & conv_std_logic_vector(-6, WEIGHT_WIDTH) & conv_std_logic_vector(11, WEIGHT_WIDTH) & conv_std_logic_vector(-5, WEIGHT_WIDTH) & conv_std_logic_vector(-12, WEIGHT_WIDTH) & conv_std_logic_vector(-4, WEIGHT_WIDTH) & conv_std_logic_vector(5, WEIGHT_WIDTH) & conv_std_logic_vector(4, WEIGHT_WIDTH) & conv_std_logic_vector(8, WEIGHT_WIDTH) & conv_std_logic_vector(4, WEIGHT_WIDTH) & conv_std_logic_vector(2, WEIGHT_WIDTH) & conv_std_logic_vector(-10, WEIGHT_WIDTH) & conv_std_logic_vector(-2, WEIGHT_WIDTH) & conv_std_logic_vector(13, WEIGHT_WIDTH) & conv_std_logic_vector(14, WEIGHT_WIDTH) & conv_std_logic_vector(-10, WEIGHT_WIDTH) & conv_std_logic_vector(9, WEIGHT_WIDTH) & conv_std_logic_vector(6, WEIGHT_WIDTH) & conv_std_logic_vector(-3, WEIGHT_WIDTH) & conv_std_logic_vector(-4, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(15, WEIGHT_WIDTH) & conv_std_logic_vector(-15, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(1, WEIGHT_WIDTH) & conv_std_logic_vector(12, WEIGHT_WIDTH) & conv_std_logic_vector(3, WEIGHT_WIDTH) & conv_std_logic_vector(-11, WEIGHT_WIDTH) & conv_std_logic_vector(-9, WEIGHT_WIDTH) & conv_std_logic_vector(11, WEIGHT_WIDTH) & conv_std_logic_vector(8, WEIGHT_WIDTH) & conv_std_logic_vector(8, WEIGHT_WIDTH) & conv_std_logic_vector(2, WEIGHT_WIDTH) & conv_std_logic_vector(14, WEIGHT_WIDTH) & conv_std_logic_vector(-6, WEIGHT_WIDTH) & conv_std_logic_vector(-7, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(19, WEIGHT_WIDTH) & conv_std_logic_vector(23, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(2, WEIGHT_WIDTH) & conv_std_logic_vector(-22, WEIGHT_WIDTH) & conv_std_logic_vector(1, WEIGHT_WIDTH) & conv_std_logic_vector(-5, WEIGHT_WIDTH) & conv_std_logic_vector(3, WEIGHT_WIDTH) & conv_std_logic_vector(3, WEIGHT_WIDTH) & conv_std_logic_vector(3, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(15, WEIGHT_WIDTH) & conv_std_logic_vector(-17, WEIGHT_WIDTH) & conv_std_logic_vector(1, WEIGHT_WIDTH) & conv_std_logic_vector(12, WEIGHT_WIDTH) & conv_std_logic_vector(-4, WEIGHT_WIDTH) & conv_std_logic_vector(3, WEIGHT_WIDTH) & conv_std_logic_vector(-5, WEIGHT_WIDTH) & conv_std_logic_vector(1, WEIGHT_WIDTH) & conv_std_logic_vector(-5, WEIGHT_WIDTH) & conv_std_logic_vector(3, WEIGHT_WIDTH) & conv_std_logic_vector(-3, WEIGHT_WIDTH) & conv_std_logic_vector(7, WEIGHT_WIDTH) & conv_std_logic_vector(25, WEIGHT_WIDTH) & conv_std_logic_vector(-14, WEIGHT_WIDTH) & conv_std_logic_vector(7, WEIGHT_WIDTH) & conv_std_logic_vector(4, WEIGHT_WIDTH) & conv_std_logic_vector(-6, WEIGHT_WIDTH) & conv_std_logic_vector(-4, WEIGHT_WIDTH) & conv_std_logic_vector(-14, WEIGHT_WIDTH) & conv_std_logic_vector(-7, WEIGHT_WIDTH) & conv_std_logic_vector(5, WEIGHT_WIDTH) & conv_std_logic_vector(-9, WEIGHT_WIDTH) & conv_std_logic_vector(6, WEIGHT_WIDTH) & conv_std_logic_vector(-2, WEIGHT_WIDTH) & conv_std_logic_vector(-4, WEIGHT_WIDTH) & conv_std_logic_vector(25, WEIGHT_WIDTH) & conv_std_logic_vector(5, WEIGHT_WIDTH) & conv_std_logic_vector(-4, WEIGHT_WIDTH) & conv_std_logic_vector(6, WEIGHT_WIDTH) & conv_std_logic_vector(14, WEIGHT_WIDTH) & conv_std_logic_vector(11, WEIGHT_WIDTH) & conv_std_logic_vector(-4, WEIGHT_WIDTH) & conv_std_logic_vector(3, WEIGHT_WIDTH) & conv_std_logic_vector(7, WEIGHT_WIDTH) & conv_std_logic_vector(2, WEIGHT_WIDTH) & conv_std_logic_vector(1, WEIGHT_WIDTH) & conv_std_logic_vector(9, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(9, WEIGHT_WIDTH) & conv_std_logic_vector(5, WEIGHT_WIDTH) & conv_std_logic_vector(5, WEIGHT_WIDTH) & conv_std_logic_vector(8, WEIGHT_WIDTH) & conv_std_logic_vector(14, WEIGHT_WIDTH) & conv_std_logic_vector(8, WEIGHT_WIDTH) & conv_std_logic_vector(-8, WEIGHT_WIDTH) & conv_std_logic_vector(16, WEIGHT_WIDTH) & conv_std_logic_vector(-4, WEIGHT_WIDTH) & conv_std_logic_vector(2, WEIGHT_WIDTH) & conv_std_logic_vector(-8, WEIGHT_WIDTH) & conv_std_logic_vector(-7, WEIGHT_WIDTH) & conv_std_logic_vector(2, WEIGHT_WIDTH) & conv_std_logic_vector(-8, WEIGHT_WIDTH) & conv_std_logic_vector(1, WEIGHT_WIDTH) & conv_std_logic_vector(10, WEIGHT_WIDTH) & conv_std_logic_vector(22, WEIGHT_WIDTH) & conv_std_logic_vector(-10, WEIGHT_WIDTH) & conv_std_logic_vector(11, WEIGHT_WIDTH) & conv_std_logic_vector(-22, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(-8, WEIGHT_WIDTH) & conv_std_logic_vector(1, WEIGHT_WIDTH) & conv_std_logic_vector(7, WEIGHT_WIDTH) & conv_std_logic_vector(-28, WEIGHT_WIDTH) & conv_std_logic_vector(3, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(1, WEIGHT_WIDTH) & conv_std_logic_vector(-9, WEIGHT_WIDTH) & conv_std_logic_vector(-1, WEIGHT_WIDTH) & conv_std_logic_vector(-15, WEIGHT_WIDTH) & conv_std_logic_vector(8, WEIGHT_WIDTH) & conv_std_logic_vector(-12, WEIGHT_WIDTH) & conv_std_logic_vector(15, WEIGHT_WIDTH) & conv_std_logic_vector(-4, WEIGHT_WIDTH) & conv_std_logic_vector(-2, WEIGHT_WIDTH) & conv_std_logic_vector(13, WEIGHT_WIDTH) & conv_std_logic_vector(23, WEIGHT_WIDTH) & conv_std_logic_vector(-10, WEIGHT_WIDTH) & conv_std_logic_vector(10, WEIGHT_WIDTH) & conv_std_logic_vector(2, WEIGHT_WIDTH) & conv_std_logic_vector(-6, WEIGHT_WIDTH) & conv_std_logic_vector(-8, WEIGHT_WIDTH) & conv_std_logic_vector(6, WEIGHT_WIDTH) & conv_std_logic_vector(3, WEIGHT_WIDTH) & conv_std_logic_vector(9, WEIGHT_WIDTH) & conv_std_logic_vector(22, WEIGHT_WIDTH) & conv_std_logic_vector(-6, WEIGHT_WIDTH),
conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH),
conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH),
conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH),
conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH) & conv_std_logic_vector(-26, WEIGHT_WIDTH),
conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH) & conv_std_logic_vector(0, WEIGHT_WIDTH)
);

end mem_settings_package;
package body mem_settings_package is
end mem_settings_package;
