library ieee;
use ieee.std_logic_1164.all;
use work.utility_package.all;
package settings_package is
constant NR_SYN                   : integer := 1;
-- decay = 2^(WEIGHT_WIDTH-1)*dt/tau
constant DECAY                    : integer_array(NR_SYN downto 0) := (15,20);

constant NR_NEURONS         : integer := 200;
constant NR_INPUT_NODES     : integer := 77;
constant CONN_FROM          : integer_matrix := ((8,24,31,92,124,155,162,163,-13,-27,-45,-75),
 (8,20,40,42,52,105,130,160,-2,-5,-23,-33),
 (9,37,101,105,126,134,191,193,-36,-53,-54,-66),
 (33,57,89,113,126,128,171,196,-11,-17,-51,-57),
 (7,25,89,91,117,133,141,180,-6,-17,-32,-40),
 (23,26,70,111,124,144,161,187,-12,-24,-28,-47),
 (19,24,72,81,84,142,156,176,-20,-24,-43,-68),
 (47,78,104,109,122,134,151,173,-29,-50,-65,-69),
 (2,84,102,105,124,131,173,190,-16,-40,-42,-69),
 (34,45,83,132,146,162,174,178,-3,-13,-19,-36),
 (25,29,61,101,112,133,141,185,-21,-67,-68,-74),
 (29,95,130,134,140,153,154,162,-15,-32,-65,-71),
 (2,31,76,89,133,165,182,194,-8,-14,-45,-67),
 (42,43,115,122,139,140,178,193,-18,-20,-47,-76),
 (5,12,15,37,163,188,193,195,-10,-31,-75,-76),
 (26,29,36,46,160,163,195,199,-1,-38,-59,-66),
 (4,54,65,86,101,131,155,183,-8,-43,-52,-76),
 (4,21,46,93,103,181,185,198,-11,-41,-62,-63),
 (47,51,88,92,124,126,127,186,-13,-37,-50,-70),
 (8,21,49,50,70,75,110,156,-13,-45,-48,-51),
 (43,44,50,72,73,138,191,198,-21,-57,-61,-73),
 (32,76,111,124,132,143,159,165,-36,-45,-61,-77),
 (19,35,36,112,154,157,164,167,-10,-52,-69,-75),
 (60,72,96,100,144,149,161,181,-35,-41,-67,-74),
 (31,56,81,101,139,152,191,194,-2,-7,-29,-51),
 (63,68,96,101,111,123,143,166,-12,-26,-41,-67),
 (12,28,32,33,46,75,195,196,-35,-39,-45,-70),
 (12,18,31,42,58,64,66,88,-39,-46,-63,-64),
 (15,46,57,62,91,105,107,114,-5,-6,-24,-41),
 (7,24,59,69,101,134,139,167,-8,-18,-21,-46),
 (3,11,46,86,91,99,181,187,-11,-20,-21,-39),
 (5,34,74,87,108,116,137,146,-17,-31,-61,-66),
 (31,56,71,83,87,116,125,186,-31,-51,-58,-70),
 (19,59,107,119,142,144,166,174,-1,-3,-6,-28),
 (4,13,33,92,111,151,154,164,-14,-15,-43,-73),
 (33,49,55,119,127,173,175,180,-8,-39,-74,-77),
 (28,37,66,93,148,159,183,192,-13,-36,-51,-56),
 (3,19,24,85,120,138,143,161,-7,-33,-47,-75),
 (16,41,45,89,121,122,135,146,-26,-35,-62,-67),
 (4,13,77,106,109,131,135,189,-33,-53,-62,-67),
 (21,22,24,30,40,93,104,152,-25,-34,-44,-64),
 (64,116,135,157,164,183,197,198,-1,-22,-24,-38),
 (10,47,55,69,81,97,175,195,-46,-61,-63,-73),
 (8,115,118,168,176,187,191,195,-3,-26,-58,-72),
 (3,107,118,121,172,174,179,183,-19,-51,-54,-62),
 (28,57,96,102,133,144,154,164,-2,-40,-51,-67),
 (18,47,66,83,85,150,183,188,-31,-53,-63,-72),
 (27,28,91,102,106,110,141,199,-19,-28,-38,-62),
 (14,55,97,107,108,122,131,160,-1,-32,-37,-52),
 (38,44,49,100,128,163,170,173,-4,-16,-56,-65),
 (1,37,39,62,78,79,132,176,-21,-25,-27,-42),
 (5,32,131,139,146,158,161,177,-2,-35,-59,-74),
 (7,10,18,41,89,106,145,181,-9,-31,-60,-62),
 (41,73,75,103,128,143,187,194,-9,-21,-71,-77),
 (3,18,30,77,109,159,164,194,-2,-5,-14,-62),
 (6,18,51,60,86,134,175,193,-5,-10,-32,-64),
 (32,43,72,86,108,117,145,178,-4,-25,-39,-68),
 (4,44,54,115,118,119,122,196,-8,-24,-28,-40),
 (12,42,78,90,115,129,142,197,-2,-7,-12,-31),
 (32,69,80,93,108,146,158,197,-20,-21,-52,-54),
 (3,10,12,57,68,82,101,180,-45,-58,-68,-72),
 (4,43,62,81,116,125,153,197,-26,-27,-36,-72),
 (117,126,149,155,164,169,174,176,-24,-45,-48,-73),
 (7,13,18,23,50,51,100,141,-29,-42,-51,-60),
 (3,6,21,33,35,105,135,137,-3,-18,-26,-44),
 (62,64,79,83,91,121,186,199,-10,-33,-42,-47),
 (15,21,62,70,82,105,168,188,-23,-37,-58,-67),
 (45,64,124,148,152,164,183,198,-1,-13,-56,-60),
 (5,10,42,69,77,119,145,190,-15,-26,-55,-70),
 (1,19,30,85,89,133,149,167,-5,-6,-14,-31),
 (60,93,104,112,136,145,166,170,-1,-39,-41,-69),
 (8,13,14,37,121,173,180,198,-6,-14,-27,-45),
 (8,29,58,74,129,135,161,189,-22,-41,-42,-63),
 (29,49,57,89,101,120,143,170,-10,-20,-37,-65),
 (9,41,67,79,81,92,136,162,-28,-30,-50,-57),
 (7,23,32,62,71,92,140,178,-26,-31,-42,-67),
 (9,11,62,107,108,137,151,199,-8,-12,-57,-63),
 (17,47,93,95,101,106,165,187,-7,-24,-48,-52),
 (3,9,32,83,126,132,138,139,-6,-12,-50,-67),
 (10,54,75,85,87,123,148,185,-14,-24,-49,-53),
 (1,49,77,88,145,163,179,189,-22,-33,-52,-66),
 (27,49,96,106,117,142,170,174,-12,-18,-60,-69),
 (4,15,33,78,91,107,125,159,-34,-35,-53,-57),
 (88,104,118,164,170,175,183,194,-28,-29,-31,-33),
 (22,27,55,63,99,143,147,161,-8,-9,-32,-33),
 (13,29,77,123,140,148,151,187,-10,-30,-34,-43),
 (7,38,55,59,70,75,76,127,-14,-18,-73,-76),
 (20,35,43,62,104,159,161,169,-4,-44,-62,-65),
 (17,23,38,48,105,124,155,173,-6,-10,-70,-74),
 (4,26,81,85,140,146,158,184,-3,-16,-25,-26),
 (34,48,52,66,67,95,105,172,-48,-63,-72,-75),
 (5,36,41,115,125,151,165,177,-37,-43,-54,-55),
 (28,54,107,122,134,142,189,190,-3,-13,-29,-55),
 (3,46,65,78,100,153,166,184,-6,-34,-55,-62),
 (1,22,34,77,81,82,131,132,-15,-21,-69,-77),
 (28,64,112,122,125,178,191,197,-1,-25,-52,-71),
 (48,111,130,149,155,181,184,200,-12,-15,-44,-75),
 (18,24,41,49,78,103,168,193,-24,-62,-68,-70),
 (3,16,54,60,84,98,113,125,-6,-21,-33,-48),
 (19,46,47,90,106,134,168,199,-2,-11,-53,-64),
 (33,35,56,64,73,125,171,191,-13,-15,-23,-43),
 (102,106,114,124,128,130,131,144,-4,-11,-17,-22),
 (49,50,59,79,145,154,169,198,-23,-55,-62,-70),
 (2,25,32,44,55,57,100,137,-7,-33,-45,-67),
 (19,50,93,102,103,112,140,172,-20,-69,-73,-77),
 (21,55,100,177,187,188,190,196,-14,-20,-22,-68),
 (6,7,43,56,59,78,150,167,-5,-15,-16,-41),
 (25,36,49,74,97,131,135,138,-37,-51,-53,-58),
 (12,41,47,48,71,73,122,145,-9,-33,-52,-59),
 (22,40,42,78,96,147,149,163,-21,-22,-71,-74),
 (38,47,54,62,105,110,152,187,-18,-20,-53,-77),
 (10,28,33,36,65,73,141,167,-42,-51,-55,-63),
 (2,40,65,83,97,138,179,185,-34,-37,-54,-67),
 (1,18,76,129,130,172,175,183,-10,-18,-35,-50),
 (11,14,65,70,111,127,159,178,-4,-16,-74,-76),
 (8,63,95,113,117,125,169,173,-16,-34,-47,-68),
 (16,53,75,124,130,140,144,184,-12,-33,-59,-61),
 (36,61,109,110,146,164,177,198,-14,-30,-63,-75),
 (1,18,70,80,95,107,117,195,-21,-31,-37,-50),
 (32,56,96,153,168,178,180,192,-2,-12,-30,-54),
 (17,20,23,40,56,108,143,177,-16,-24,-44,-55),
 (27,41,46,95,106,161,167,184,-9,-24,-34,-65),
 (19,57,132,136,139,161,192,194,-11,-35,-46,-77),
 (19,20,81,115,122,167,182,199,-2,-11,-39,-76),
 (23,39,40,82,119,127,143,170,-34,-36,-50,-55),
 (13,44,101,118,142,160,162,171,-13,-39,-46,-48),
 (5,6,23,65,72,78,103,172,-14,-30,-40,-46),
 (29,77,79,82,84,104,167,179,-36,-42,-55,-58),
 (63,89,99,103,129,146,160,163,-18,-25,-70,-73),
 (4,20,79,101,135,145,175,185,-19,-27,-34,-46),
 (10,15,16,22,36,49,102,138,-2,-22,-51,-76),
 (31,40,104,115,127,154,185,196,-24,-52,-56,-60),
 (43,92,101,115,131,172,178,197,-7,-9,-37,-46),
 (18,33,75,90,103,108,121,148,-18,-23,-61,-63),
 (2,4,21,24,31,87,109,134,-8,-47,-53,-70),
 (31,85,105,126,129,146,148,171,-4,-9,-31,-70),
 (3,24,34,35,119,122,177,196,-7,-14,-23,-30),
 (47,69,109,140,153,168,174,180,-9,-14,-52,-77),
 (53,54,56,62,94,115,164,173,-7,-18,-25,-60),
 (7,31,35,71,137,143,145,157,-17,-35,-36,-61),
 (15,20,25,47,53,56,150,169,-8,-35,-40,-56),
 (1,14,41,75,93,100,190,197,-6,-19,-24,-43),
 (42,75,89,113,159,160,169,196,-24,-25,-50,-74),
 (38,52,54,112,116,129,164,184,-7,-17,-26,-61),
 (1,52,60,61,81,97,117,174,-28,-33,-65,-70),
 (54,75,117,123,148,179,180,189,-4,-25,-34,-45),
 (9,15,25,41,64,75,94,105,-42,-46,-68,-76),
 (2,3,10,35,57,96,101,199,-27,-44,-61,-64),
 (111,124,126,133,138,160,162,197,-12,-16,-56,-68),
 (47,95,121,127,149,182,186,200,-8,-27,-63,-65),
 (8,11,38,44,98,139,143,167,-50,-52,-57,-58),
 (7,12,34,71,99,117,162,185,-8,-15,-46,-70),
 (9,51,58,102,105,107,124,196,-45,-47,-69,-71),
 (1,29,36,73,77,165,180,193,-12,-21,-53,-64),
 (9,34,39,119,154,197,198,199,-2,-5,-14,-20),
 (31,61,83,131,174,178,181,195,-1,-4,-9,-71),
 (46,48,63,75,78,80,85,139,-16,-37,-53,-73),
 (23,27,30,34,60,76,103,145,-23,-43,-46,-59),
 (3,21,29,41,56,96,138,177,-13,-31,-36,-69),
 (41,56,68,122,143,183,186,199,-15,-36,-72,-74),
 (20,43,65,112,123,156,177,193,-10,-11,-21,-42),
 (75,91,97,101,102,139,142,159,-16,-66,-68,-75),
 (45,47,96,127,133,138,146,199,-9,-47,-57,-63),
 (1,29,67,98,104,153,173,184,-1,-43,-50,-67),
 (2,46,90,108,113,127,146,177,-16,-47,-66,-77),
 (37,43,47,56,81,97,104,128,-10,-38,-46,-63),
 (8,13,48,84,95,124,196,198,-7,-13,-48,-55),
 (7,35,40,64,134,136,139,162,-18,-45,-56,-61),
 (16,31,33,58,90,126,154,173,-29,-35,-36,-52),
 (19,40,45,53,95,124,143,169,-2,-16,-27,-53),
 (4,27,30,34,35,128,184,189,-11,-14,-34,-41),
 (12,19,31,41,52,112,129,167,-12,-48,-69,-73),
 (15,20,56,75,114,126,178,180,-3,-13,-52,-67),
 (4,25,35,48,64,88,152,161,-22,-38,-53,-65),
 (69,84,96,143,162,177,180,182,-53,-69,-70,-76),
 (25,46,82,86,105,130,144,165,-9,-42,-64,-72),
 (7,9,20,42,76,147,149,192,-21,-26,-71,-77),
 (3,25,90,101,111,120,161,195,-15,-27,-40,-73),
 (68,69,73,122,127,132,138,195,-2,-4,-58,-68),
 (2,9,15,39,78,142,145,180,-13,-15,-46,-57),
 (27,111,119,133,171,179,187,197,-12,-35,-36,-71),
 (11,58,68,80,94,146,182,197,-5,-29,-45,-48),
 (26,33,42,55,83,99,100,188,-4,-20,-33,-75),
 (5,38,59,67,82,125,172,182,-15,-37,-54,-69),
 (14,33,90,106,136,148,170,190,-21,-40,-59,-73),
 (3,14,15,76,118,157,166,174,-47,-53,-71,-73),
 (34,65,96,133,137,144,165,179,-7,-12,-25,-75),
 (55,56,88,93,97,147,157,200,-7,-13,-25,-71),
 (26,32,51,97,108,175,187,200,-16,-24,-40,-54),
 (62,78,95,113,117,118,176,180,-7,-36,-46,-64),
 (32,40,53,73,99,113,165,168,-13,-22,-51,-69),
 (71,78,84,157,159,178,183,184,-10,-11,-36,-61),
 (24,38,59,62,98,126,130,178,-9,-15,-49,-75),
 (69,82,113,120,122,178,196,200,-36,-40,-65,-75),
 (6,68,133,152,180,189,197,199,-4,-34,-43,-69),
 (34,68,69,83,93,119,123,139,-6,-26,-45,-46),
 (13,51,77,83,123,166,183,199,-5,-39,-40,-75),
 (5,30,47,101,102,121,158,180,-17,-34,-67,-69),
 (11,17,18,61,136,151,164,193,-8,-24,-65,-76),
 (14,22,63,122,131,136,145,146,-8,-14,-26,-36));
 constant NR_OUTPUT_NODES    : integer := 200;
constant OUTPUT_NODES       : integer_array := (1,2,3,4,5,6,7,8,9,10,11,12,13,14,15,16,17,18,19,20,21,22,23,24,25,26,27,28,29,30,31,32,33,34,35,36,37,38,39,40,41,42,43,44,45,46,47,48,49,50,51,52,53,54,55,56,57,58,59,60,61,62,63,64,65,66,67,68,69,70,71,72,73,74,75,76,77,78,79,80,81,82,83,84,85,86,87,88,89,90,91,92,93,94,95,96,97,98,99,100,101,102,103,104,105,106,107,108,109,110,111,112,113,114,115,116,117,118,119,120,121,122,123,124,125,126,127,128,129,130,131,132,133,134,135,136,137,138,139,140,141,142,143,144,145,146,147,148,149,150,151,152,153,154,155,156,157,158,159,160,161,162,163,164,165,166,167,168,169,170,171,172,173,174,175,176,177,178,179,180,181,182,183,184,185,186,187,188,189,190,191,192,193,194,195,196,197,198,199,200);
 constant SYNAPSE_MAP        : integer_matrix := ((0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12),
 (0,12));
 end settings_package;
package body settings_package is
end settings_package;
