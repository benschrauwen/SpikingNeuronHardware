library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_signed.all;
use work.settings_package.all;
package intercon_mem_package is
constant intercon_mem : con_mem_type := (
"10000111011",
"10000100000",
"10000011110",
"10000110001",
"10000100010",
"10000110101",
"10000001100",
"10001001011",
"10000111001",
"10000110011",
"10001001011",
"10001001000",
"10001000001",
"10001001010",
"10001010001",
"10000111110",
"10001001001",
"10000101100",
"10001001101",
"10001001001",
"10000110001",
"10001001001",
"10001001011",
"10000101101",
"10000010011",
"10001000110",
"10001001110",
"10001010000",
"10001001000",
"10001000100",
"10000111110",
"10001001000",
"10001001010",
"10000011110",
"10000110100",
"10001010000",
"10001001101",
"10001000110",
"10000100110",
"10001010010",
"10001000000",
"10000111111",
"10000101010",
"10000111100",
"10000110000",
"10000100001",
"10000100111",
"10001001110",
"10000001001",
"10000100101",
"10000111011",
"10000110010",
"10000101101",
"10001010000",
"10000111100",
"10000001100",
"10001000100",
"10000110011",
"10000110101",
"10001000110",
"10000110101",
"10000110001",
"10001001110",
"10001010010",
"10001000110",
"10000100110",
"10001000011",
"10001001111",
"10000110110",
"10000111110",
"10001000100",
"10000101000",
"10001000110",
"10001000111",
"10000110001",
"10000110100",
"10000111101",
"10000011111",
"10000111000",
"10001000101",
"10000111101",
"10001001000",
"10001001010",
"10000101011",
"10000110100",
"10000111001",
"10001000001",
"10000011111",
"10000111111",
"10001001001",
"10001010010",
"10001001100",
"10001000010",
"10000111110",
"10001001110",
"10000110111",
"10000110111",
"10000010010",
"10000101001",
"10000011000",

"10000010100",
"10000011100",
"10000000111",
"10000000101",
"10000001011",
"10000100001",
"10000001001",
"10000001011",
"10000101110",
"10000110001",
"10000000101",
"10000100100",
"10000101000",
"10000101011",
"10000010100",
"10000101010",
"10000000110",
"10000100100",
"10000111011",
"10000101010",
"10000101101",
"10000010110",
"10000011110",
"10000100101",
"10000001001",
"10000110100",
"10001001011",
"10000011000",
"10000100101",
"10000111011",
"10000101101",
"10000101100",
"10000110100",
"10000001111",
"10000010000",
"10001001011",
"10000101000",
"10000001010",
"10000100101",
"10000011101",
"10000000101",
"10000011001",
"10000011101",
"10000001101",
"10000001100",
"10000011100",
"10000011000",
"10001001000",
"10000000111",
"10000011100",
"10000100101",
"10000001100",
"10000101011",
"10000101110",
"10000110000",
"10000001010",
"10000101011",
"10000100101",
"10000101000",
"10000101100",
"10000101001",
"10000100001",
"10000111010",
"10001000110",
"10000110010",
"10000011110",
"10000101000",
"10001001000",
"10000000101",
"10000100010",
"10000111000",
"10000100011",
"10000110010",
"10000000111",
"10000110000",
"10000100011",
"10000110111",
"10000011010",
"10000001111",
"10001000010",
"10000110110",
"10000011011",
"10000011101",
"10000100111",
"10000010110",
"10000001011",
"10000010000",
"10000001010",
"10000100100",
"10000010011",
"10000111011",
"10000111000",
"10000110111",
"10000010101",
"10000100010",
"10000010101",
"10000110110",
"10000001001",
"10000100011",
"10000000110",

"01000110101",
"01001001000",
"01001011010",
"01000101010",
"01000111011",
"01000001100",
"01000010101",
"01000110111",
"01001100001",
"01001011111",
"01001011011",
"00110110011",
"00110101111",
"01001100011",
"01001011111",
"01000111110",
"01000001101",
"01001011000",
"01001011110",
"01000000001",
"01000111000",
"01000111111",
"01000011101",
"01000110101",
"01001000100",
"01001001100",
"01001011010",
"01001100000",
"01001100010",
"01001011100",
"01000001100",
"01000100000",
"01001010101",
"00111010110",
"01000111101",
"01000010011",
"01000101101",
"01001100001",
"01000000111",
"01001011000",
"01000100010",
"00100101111",
"00110110101",
"01001011011",
"01001010000",
"01000100101",
"01001011100",
"01001001110",
"01000110110",
"01001000101",
"01001011111",
"01001010110",
"01001100011",
"01000110110",
"01001000001",
"01000111000",
"01000010001",
"01001011111",
"01001011011",
"01001010010",
"01000001110",
"01001100000",
"01001010111",
"01001001001",
"01001010100",
"00111100010",
"00111100011",
"01000111101",
"01001000001",
"01001001101",
"01000010100",
"01000111011",
"01000101110",
"01000111011",
"01000111101",
"01001010010",
"01000100001",
"00111010010",
"01001100010",
"01001010010",
"01000000110",
"01001000100",
"01001011110",
"01000101101",
"00111010011",
"01001011101",
"01000111000",
"01000100100",
"01001011000",
"01000100100",
"00111011001",
"00110001000",
"01001000000",
"00110111110",
"01000101111",
"01001001100",
"01001010110",
"01000110101",
"01001001011",
"00110001101",

"00110011110",
"00110100100",
"01000101011",
"01000100000",
"01000110111",
"00111001101",
"01000000111",
"01000010110",
"01001000111",
"01000111001",
"00101010111",
"00110010110",
"00110000101",
"01001000001",
"01001000111",
"00111000001",
"01000001000",
"01000101111",
"00110111010",
"00111010001",
"00111011100",
"01000010100",
"00110101010",
"01000010111",
"01001000011",
"01001000001",
"01000111001",
"01001011111",
"01000100001",
"00110111111",
"01000001010",
"00110010100",
"00111001001",
"00110110111",
"01000101110",
"00110001111",
"01000011000",
"01001000011",
"00111000010",
"01000000001",
"01000010110",
"00011010000",
"00110100000",
"01001010001",
"01001001110",
"01000100011",
"01000010101",
"01000110010",
"01000110100",
"00110101111",
"00111001011",
"00111011111",
"00110111001",
"01000100111",
"01000101010",
"00111000011",
"00111000000",
"01001010010",
"00111010111",
"01001001010",
"00111010100",
"01001011101",
"01000111001",
"01000111011",
"01000101110",
"00111000001",
"00111010110",
"01000110001",
"01000101011",
"01001001000",
"01000000001",
"00111001101",
"00111011101",
"00111000110",
"01000000011",
"00111011110",
"00101011001",
"00110111111",
"01001001111",
"01000010100",
"00110000010",
"01001000001",
"01000010110",
"01000010100",
"00110100011",
"01001010000",
"01000011010",
"01000001101",
"01001010100",
"01000010011",
"00111001010",
"00101010010",
"01000110001",
"00110100111",
"01000000000",
"01000100100",
"01001010001",
"00111100010",
"00101001011",
"00101001111",

"00101011001",
"00100100011",
"00111010111",
"01000001111",
"01000100010",
"00110100110",
"01000000101",
"00110111001",
"01000000001",
"01000111000",
"00100011010",
"00110001101",
"00100101001",
"01000011101",
"01000101010",
"00100110011",
"00110100111",
"01000000000",
"00110101000",
"00110111111",
"00110100010",
"01000010001",
"00100110100",
"00111010010",
"01000111110",
"01000010111",
"00111001101",
"01001001110",
"01000001110",
"00100111101",
"01000000111",
"00110000001",
"00110100100",
"00110010110",
"01000011111",
"00110000111",
"01000001010",
"00111010101",
"00110010111",
"00110001110",
"00110100010",
"00010101011",
"00101011101",
"00110100011",
"01001000110",
"01000100010",
"00110001011",
"01000011110",
"01000101001",
"00101000101",
"00110111100",
"00111010000",
"00110001110",
"01000100101",
"01000100100",
"00110101110",
"00100011111",
"01001001111",
"00110000000",
"01000110000",
"00110101011",
"01001011000",
"01000110000",
"01000110000",
"01000001101",
"00110101011",
"00110110011",
"01000100001",
"00111011011",
"01000010101",
"00101100010",
"00110001111",
"00111001001",
"00110100101",
"00111010000",
"00111001111",
"00100010110",
"00110100101",
"00111000001",
"01000010000",
"00100111110",
"00110110011",
"00110101110",
"01000000110",
"00110011101",
"01000111011",
"00111000111",
"00111010110",
"01000101011",
"01000001010",
"00100001111",
"00100101110",
"01000000111",
"00110001100",
"00100111010",
"00111010101",
"00111001100",
"00110111110",
"00101000011",
"00100111101",

"00101000100",
"00100001111",
"00111000000",
"00110111011",
"01000000001",
"00110011010",
"00110110001",
"00110101011",
"00110011100",
"01000000100",
"00100010111",
"00100110011",
"00100010100",
"00110111101",
"00110100001",
"00011011111",
"00110100101",
"00101011111",
"00101001010",
"00110101110",
"00101001010",
"01000000011",
"00100100111",
"00110110001",
"00110001110",
"00111100001",
"00110111000",
"01000101111",
"00110101111",
"00011000101",
"00111001001",
"00100110001",
"00110001011",
"00100110110",
"01000000111",
"00110000110",
"00110100111",
"00111000001",
"00100001100",
"00100101101",
"00110010110",
"00010001001",
"00100101010",
"00110000010",
"00101000001",
"00110111111",
"00100101001",
"01000010111",
"01000001110",
"00100101101",
"00101100011",
"00110001000",
"00101100001",
"01000000000",
"00110111100",
"00101001001",
"00100001100",
"00111011111",
"00101011101",
"00110111101",
"00110011101",
"00111001011",
"01000100110",
"00111000010",
"01000000111",
"00110000100",
"00110001011",
"01000001100",
"00110000001",
"00110101001",
"00101011000",
"00101001110",
"00101010100",
"00100111000",
"00111001011",
"00110111101",
"00100010010",
"00101000010",
"00100110101",
"01000000111",
"00100100110",
"00011010101",
"00110101011",
"00111100001",
"00101100011",
"00111010101",
"00110011010",
"00111000010",
"01000000001",
"00110111110",
"00011011110",
"00010100011",
"01000000100",
"00101001010",
"00100110000",
"00110011111",
"00101010010",
"00101010111",
"00100111101",
"00100110000",

"00100100010",
"00011100001",
"00110101100",
"00110010100",
"00111100011",
"00100010101",
"00110100001",
"00101000001",
"00101011011",
"00101011101",
"00011100010",
"00011001101",
"00100000010",
"00110100000",
"00100111010",
"00010011001",
"00110010111",
"00100101110",
"00100010100",
"00110010001",
"00100110100",
"00110111011",
"00100010111",
"00110100111",
"00110000111",
"00111000101",
"00110001010",
"00111011110",
"00100000001",
"00010111111",
"00110011010",
"00010010001",
"00100111100",
"00011000101",
"00110101011",
"00101100011",
"00101011011",
"00110011001",
"00001010000",
"00100101011",
"00100110111",
"00001011110",
"00100001011",
"00011100001",
"00100000110",
"00101011011",
"00011011101",
"00101000000",
"01000000111",
"00011011000",
"00101010101",
"00100111101",
"00010011001",
"00101011010",
"00110111001",
"00101000101",
"00011011111",
"00111011101",
"00101001110",
"00101100011",
"00110010100",
"00110010110",
"00110101000",
"00110111101",
"00111010010",
"00100101000",
"00010110110",
"01000001000",
"00100111111",
"00110000101",
"00100100111",
"00011011111",
"00100110111",
"00100010000",
"00100011001",
"00100110101",
"00100000101",
"00100100111",
"00100001110",
"00110010100",
"00100100001",
"00010101100",
"00110101010",
"00111010100",
"00101000010",
"00110000010",
"00101100000",
"00110110010",
"00110010001",
"00110100100",
"00010110110",
"00000111011",
"00100101001",
"00101000110",
"00100101011",
"00101010001",
"00100011100",
"00101000011",
"00100001000",
"00100101001",

"00011000001",
"00010111111",
"00010101101",
"00100110100",
"00010110110",
"00100000001",
"00110000101",
"00011001111",
"00101001100",
"00101011001",
"00011001100",
"00001001101",
"00010110010",
"00110001111",
"00011000001",
"00001100010",
"00101010010",
"00011011001",
"00100000011",
"00100101111",
"00011011100",
"00110101101",
"00010000100",
"00110100100",
"00011011101",
"00110000011",
"00110001001",
"00010101000",
"00011010010",
"00010011010",
"00100100111",
"00010010000",
"00100000010",
"00010111111",
"00101011010",
"00100101010",
"00101000000",
"00011010110",
"00000111011",
"00010110100",
"00010100101",
"00001001111",
"00011010011",
"00011001000",
"00100000001",
"00101000101",
"00011010101",
"00100110110",
"00101011100",
"00010010110",
"00101001011",
"00100101110",
"00010000111",
"00100011010",
"00110100001",
"00011011111",
"00001100000",
"00100100001",
"00101001000",
"00100110111",
"00101010101",
"00110000101",
"00101011010",
"00110001110",
"00100110101",
"00010100011",
"00001100011",
"00101000011",
"00010111100",
"00101001111",
"00010111100",
"00011001111",
"00100101110",
"00010110011",
"00010100010",
"00100001111",
"00011011111",
"00100010010",
"00011001011",
"00110001001",
"00100000010",
"00010100111",
"00011011110",
"00110100000",
"00100011101",
"00101010011",
"00011100011",
"00101100011",
"00110001010",
"00001011001",
"00010001001",
"00000101101",
"00100001111",
"00100110110",
"00100000110",
"00100111101",
"00011010011",
"00100110101",
"00011001111",
"00010001101",

"00010111111",
"00010110000",
"00010010110",
"00100000110",
"00000110001",
"00011001001",
"00100000001",
"00010101110",
"00101000110",
"00100100101",
"00010101011",
"00001000100",
"00010001000",
"00100010100",
"00010110011",
"00001001011",
"00010110001",
"00001000101",
"00010111011",
"00100001001",
"00010101101",
"00100100000",
"00001001101",
"00100100011",
"00001001001",
"00100100100",
"00101001100",
"00010010010",
"00010011100",
"00010001000",
"00011100000",
"00010001000",
"00011011111",
"00010110001",
"00101010100",
"00011001110",
"00100101111",
"00010111101",
"00000110100",
"00010101111",
"00010011001",
"00001000000",
"00010011101",
"00010110000",
"00011100010",
"00011001111",
"00011001000",
"00100000111",
"00001001011",
"00001000011",
"00101001000",
"00100000011",
"00001011111",
"00010101110",
"00011011001",
"00010111100",
"00001000001",
"00100000111",
"00100110110",
"00100110101",
"00100011101",
"00100000110",
"00100101110",
"00101000100",
"00100010000",
"00001100011",
"00000101110",
"00100011110",
"00001010001",
"00100000011",
"00010110100",
"00001010111",
"00100101101",
"00010010001",
"00010011110",
"00010011000",
"00010110011",
"00011001000",
"00011001000",
"00110000000",
"00010010110",
"00010010111",
"00010101110",
"00110000101",
"00011011000",
"00011100011",
"00010100101",
"00100000111",
"00101011111",
"00001010100",
"00010000110",
"00000101011",
"00100001101",
"00011100011",
"00011010101",
"00100101011",
"00010001100",
"00010100101",
"00010010000",
"00001011111",

"00001011100",
"00010101111",
"00001100000",
"00000111100",
"00000101011",
"00001001001",
"00010100100",
"00010011111",
"00100111011",
"00100000000",
"00010010010",
"00000111110",
"00001011001",
"00100001101",
"00001001110",
"00000110000",
"00010001100",
"00000100010",
"00010100100",
"00001011100",
"00010011011",
"00010000010",
"00000101100",
"00100011000",
"00000111001",
"00010011011",
"00100000001",
"00010001110",
"00001010001",
"00000101101",
"00011011001",
"00010000001",
"00001000111",
"00001001010",
"00101001111",
"00000110011",
"00100100110",
"00010110010",
"00000101010",
"00010010001",
"00010010010",
"00000111001",
"00010000101",
"00010001000",
"00011000000",
"00010111110",
"00010010011",
"00000110110",
"00000110000",
"00000001111",
"00101000000",
"00011010101",
"00000111010",
"00010000101",
"00010101111",
"00010110111",
"00000101101",
"00010000100",
"00010100110",
"00001010100",
"00001001011",
"00010011111",
"00011001110",
"00100010100",
"00011010010",
"00000101010",
"00000011101",
"00011100001",
"00000101010",
"00001010111",
"00001000111",
"00001000000",
"00100100111",
"00001100001",
"00010011001",
"00010010011",
"00001011100",
"00010110110",
"00001001100",
"00101001100",
"00001100011",
"00010010010",
"00010010111",
"00100110011",
"00010000101",
"00010101001",
"00010100010",
"00011000111",
"00100010000",
"00001010000",
"00010000001",
"00000011011",
"00100000010",
"00010100111",
"00010011111",
"00100100100",
"00001000101",
"00010011100",
"00010000100",
"00001001011",

"00000110111",
"00001000001",
"00001010000",
"00000000111",
"00000010110",
"00000101111",
"00010010010",
"00010000010",
"00010001011",
"00011011111",
"00000011010",
"00000111101",
"00000000110",
"00001011011",
"00000110000",
"00000101111",
"00001010110",
"00000011101",
"00010010101",
"00000110110",
"00010000011",
"00000111111",
"00000011110",
"00010101011",
"00000110001",
"00000111101",
"00010111010",
"00001001011",
"00001000100",
"00000001010",
"00010110111",
"00001100000",
"00001000000",
"00001000110",
"00100100011",
"00000101010",
"00010001001",
"00010010100",
"00000010010",
"00000110100",
"00001011110",
"00000110111",
"00001010111",
"00000010001",
"00000010111",
"00010000000",
"00010000111",
"00000110001",
"00000101111",
"00000000011",
"00100000101",
"00011010100",
"00000101101",
"00000010100",
"00000100010",
"00010100010",
"00000011011",
"00000111010",
"00010011001",
"00000110001",
"00000111111",
"00010001101",
"00010110110",
"00010101111",
"00010011011",
"00000011010",
"00000010000",
"00000010111",
"00000011001",
"00000010001",
"00000010101",
"00000110111",
"00001011110",
"00000010010",
"00001011010",
"00000100001",
"00001000001",
"00010010110",
"00000100011",
"00000110110",
"00000101101",
"00010001110",
"00001100010",
"00100011010",
"00000101100",
"00000001001",
"00010100000",
"00001011011",
"00100000010",
"00000001011",
"00000100100",
"00000001101",
"00000110011",
"00001010100",
"00010010000",
"00010101011",
"00000111011",
"00001010111",
"00001011011",
"00001001001",

"00000010101",
"00000111111",
"00000011101",
"00000000001",
"00000010010",
"00000000111",
"00000011101",
"00000001010",
"00000100100",
"00010111010",
"00000000001",
"00000101110",
"00000000100",
"00000100111",
"00000011100",
"00000101001",
"00000000001",
"00000011001",
"00000010110",
"00000000110",
"00000011000",
"00000111001",
"00000000000",
"00010000100",
"00000000101",
"00000100010",
"00010001001",
"00001000001",
"00000110110",
"00000000011",
"00001100001",
"00000001000",
"00000111001",
"00000000000",
"00010110010",
"00000011010",
"00001010101",
"00001001110",
"00000000011",
"00000110010",
"00001011000",
"00000101100",
"00001001110",
"00000001000",
"00000000000",
"00001000100",
"00000110000",
"00000010111",
"00000101110",
"00000000001",
"00011011111",
"00001011111",
"00000001101",
"00000000000",
"00000000001",
"00010000001",
"00000001100",
"00000101110",
"00010000011",
"00000110000",
"00000010010",
"00001000001",
"00000000101",
"00000001100",
"00010010000",
"00000000010",
"00000001101",
"00000010000",
"00000010001",
"00000000000",
"00000010001",
"00000110000",
"00001001000",
"00000001000",
"00001010010",
"00000010110",
"00000001111",
"00010010101",
"00000010111",
"00000000111",
"00000100100",
"00001100000",
"00000110111",
"00100001000",
"00000100101",
"00000000010",
"00001100011",
"00000100100",
"00010001000",
"00000000100",
"00000000001",
"00000000001",
"00000100010",
"00000001111",
"00010001000",
"00010100001",
"00000110101",
"00001001100",
"00000001001",
"00000010011",


"10000110001",
"10000111111",
"10000100010",
"10000101001",
"10000110110",
"10000101101",
"10000101011",
"10000011110",
"10001001101",
"10000010011",
"10000110111",
"10000111000",
"10001001010",
"10001000111",
"10001001011",
"10000011101",
"10001010000",
"10001000101",
"10000100111",
"10001010001",
"10000111000",
"10001001011",
"10000010010",
"10000111111",
"10001000100",
"10001001010",
"10000110101",
"10000011100",
"10000011100",
"10001010000",
"10001001101",
"10001000011",
"10000010011",
"10001001000",
"10001001011",
"10001010001",
"10000011101",
"10001001001",
"10001001111",
"10000111100",
"10000110111",
"10000101101",
"10001000100",
"10000100000",
"10000101011",
"10000100111",
"10000100000",
"10000100001",
"10000101110",
"10001000001",
"10000101010",
"10000110110",
"10000011010",
"10001001001",
"10000111010",
"10000100110",
"10000100001",
"10001001000",
"10000111111",
"10000111110",
"10000111010",
"10000110101",
"10000110011",
"10000111100",
"10000111100",
"10000111110",
"10000111011",
"10001001111",
"10001001101",
"10000110001",
"10001010001",
"10000100100",
"10000100010",
"10001001101",
"10001000101",
"10000111011",
"10000011111",
"10001000101",
"10001000010",
"10001001000",
"10001000101",
"10001010001",
"10000110110",
"10000111011",
"10000110100",
"10000100110",
"10000101111",
"10001001100",
"10001001011",
"10000100100",
"10000110000",
"10000011111",
"10000111111",
"10001010010",
"10000011110",
"10001000010",
"10000101011",
"10001000110",
"10001000001",
"10000011001",

"10000100111",
"10000110111",
"10000001000",
"10000101000",
"10000101000",
"10000000110",
"10000011000",
"10000010011",
"10000111010",
"10000000110",
"10000001100",
"10000000110",
"10000011110",
"10000101101",
"10000001001",
"10000001011",
"10001001011",
"10000011001",
"10000100110",
"10001001100",
"10000011011",
"10001000101",
"10000010000",
"10000110111",
"10000111000",
"10000101000",
"10000101100",
"10000000101",
"10000011010",
"10000010100",
"10000100111",
"10000010011",
"10000001110",
"10000100010",
"10000001000",
"10000000101",
"10000001110",
"10000011100",
"10000101100",
"10000010100",
"10000101011",
"10000100000",
"10000110100",
"10000011011",
"10000011000",
"10000011111",
"10000010010",
"10000011011",
"10000010100",
"10000011001",
"10000010011",
"10000001100",
"10000001110",
"10000111010",
"10000000110",
"10000011001",
"10000011100",
"10000100111",
"10000100011",
"10000110111",
"10000001110",
"10000000110",
"10000001111",
"10000000111",
"10000100000",
"10000101011",
"10000010111",
"10001001110",
"10000100110",
"10000100001",
"10000010011",
"10000000110",
"10000100001",
"10000011110",
"10000000110",
"10000100011",
"10000001010",
"10000100110",
"10000111101",
"10000110111",
"10000111100",
"10000110010",
"10000001100",
"10000101110",
"10000010011",
"10000011110",
"10000001110",
"10000011010",
"10001001000",
"10000001111",
"10000010001",
"10000000110",
"10000010010",
"10000011111",
"10000001111",
"10000010110",
"10000010000",
"10000110000",
"10000001000",
"10000001011",

"01001010010",
"01001010110",
"01001100001",
"01001001000",
"01001100001",
"01001011100",
"01000101001",
"01001010011",
"01001011101",
"01001010010",
"01000010011",
"01001001110",
"01001001011",
"01000110101",
"01001011101",
"01001000000",
"01000000010",
"01001010111",
"00111001101",
"01000000011",
"01001010110",
"01000101000",
"01000111011",
"01001010100",
"01000100011",
"00110111100",
"00111010001",
"00111011011",
"01001011000",
"01000100010",
"01001001011",
"00111010010",
"01001010101",
"01000011001",
"01001010011",
"01000101110",
"01000001110",
"01000010111",
"01001100001",
"01001011101",
"01001000110",
"01001000001",
"01001010001",
"01001100000",
"01001010101",
"01000111111",
"01000111100",
"01000110101",
"01000110111",
"01001010110",
"01001001100",
"01000110111",
"01000101110",
"01001001101",
"01001011101",
"01001100011",
"01000101111",
"01000101011",
"01001010001",
"01001001111",
"01000001111",
"01000110110",
"00111011010",
"01001000000",
"01001001001",
"01000111000",
"01001100010",
"01000110000",
"01000011110",
"01001000011",
"01000110110",
"01000101101",
"01001011000",
"01001000001",
"00110101001",
"00110110111",
"01000111111",
"01001001110",
"01000011110",
"01000100001",
"01000111000",
"01001011001",
"01000111000",
"01000110101",
"01001001001",
"00111100010",
"01000101100",
"01000011011",
"01001001110",
"01001000000",
"01001010000",
"01001001011",
"00111010011",
"01001011100",
"01001010100",
"01001010110",
"01000111110",
"01001010101",
"01001011001",
"01001010011",

"01001001101",
"01001000101",
"01001010011",
"01001000000",
"01000101011",
"01000010001",
"00110110100",
"01000110100",
"01001010101",
"01001000000",
"00111100011",
"01001000011",
"01001000011",
"00111010110",
"01001011011",
"01000110011",
"00101000101",
"01001000000",
"00100110101",
"00111011101",
"01001010100",
"01000100111",
"01000100111",
"01000100101",
"01000001110",
"00100110001",
"00110110111",
"00110010110",
"01000101111",
"00111100010",
"01000011010",
"00110101011",
"01001010100",
"01000000110",
"01000110010",
"00111010100",
"00110100110",
"01000001110",
"01000111100",
"01000000110",
"01000010010",
"01000110111",
"01000111011",
"01001011110",
"00111001010",
"00111001000",
"01000001000",
"01000110010",
"00111100010",
"01000111000",
"01000000011",
"00111000100",
"00111001100",
"01001001001",
"01000111001",
"01001000011",
"00100100011",
"01000000001",
"01000100110",
"01001001100",
"00111011010",
"01000110101",
"00110101001",
"01000000111",
"01001000000",
"00111011000",
"01000110001",
"01000100110",
"00110110001",
"01000001011",
"01000100001",
"00111001011",
"00111100011",
"00111010110",
"00110100111",
"00110101010",
"01000001000",
"01000001101",
"01000010110",
"01000010100",
"00111010111",
"01000110010",
"00110111110",
"01000101010",
"01000100111",
"00110110101",
"01000101000",
"01000000000",
"00111011110",
"01000111110",
"00111000111",
"00110110110",
"00101100000",
"01001001110",
"01001001101",
"00110111011",
"00111011101",
"00111100001",
"00101011110",
"01000001101",

"01001000000",
"00111001101",
"01001000100",
"00111000000",
"01000101010",
"01000000010",
"00110101101",
"00111001110",
"01000101001",
"00110111100",
"00111001111",
"01000011101",
"01000110100",
"00111000111",
"01001010010",
"00111000110",
"00100001100",
"01000001101",
"00010110101",
"00110011110",
"01000110111",
"00111011010",
"01000011011",
"00111011110",
"00100101100",
"00100101010",
"00110010000",
"00110010010",
"01000101101",
"00110010111",
"00110110101",
"00101100010",
"01001000101",
"00100010001",
"01000101010",
"00101001000",
"00110010100",
"00111000011",
"01000110011",
"01000000011",
"00111000001",
"01000100101",
"01000100111",
"01001011001",
"00110010010",
"00110010000",
"00111100011",
"01000000001",
"00111011111",
"01000000111",
"00101001100",
"00110010010",
"00110111011",
"01000010110",
"00110111100",
"01000101001",
"00100011011",
"00111010110",
"01000000110",
"01000110100",
"00111010010",
"01000101101",
"00110010101",
"01000000101",
"00110010000",
"00111010111",
"01000010011",
"01000000010",
"00110010100",
"00111100001",
"00111011111",
"00110001010",
"00111010000",
"00111000000",
"00110100000",
"00101001010",
"00111100001",
"00110111001",
"00100111110",
"01000000100",
"00110110111",
"01000100101",
"00110100010",
"01000000001",
"01000001110",
"00100100010",
"01000001001",
"00110010101",
"00111000010",
"01000101000",
"00110110101",
"00110000010",
"00101000101",
"01001001101",
"00111011100",
"00110100010",
"00110011010",
"00110001100",
"00100111101",
"00111100000",

"00111001000",
"00110100110",
"00100101011",
"00110100110",
"00111100011",
"00111011000",
"00110010000",
"00110100100",
"01000100101",
"00110010111",
"00110100111",
"00110000000",
"01000101000",
"00110111010",
"01000001111",
"00110101001",
"00100000010",
"00110100010",
"00010100101",
"00101011110",
"00111001000",
"00110110000",
"00101010111",
"00110011011",
"00100000001",
"00100100010",
"00101011100",
"00100000011",
"01000001001",
"00110000000",
"00110110100",
"00101010011",
"01000101101",
"00011100011",
"01000011011",
"00100110100",
"00110001111",
"00110010010",
"01000100101",
"01000000010",
"00101100000",
"00110010010",
"00101010111",
"01000100111",
"00101000000",
"00101011010",
"00111010101",
"00110001100",
"00110101001",
"00110110101",
"00100010001",
"00100010100",
"00101011000",
"00110011010",
"00110101101",
"00110111011",
"00011010001",
"00110100010",
"01000000011",
"00111001010",
"00111000111",
"00110110001",
"00110000100",
"00111011100",
"00110000110",
"00110110100",
"01000010010",
"00110010111",
"00110000111",
"00110011011",
"00101010111",
"00100101110",
"00110100101",
"00101011101",
"00110011101",
"00011100011",
"00110111100",
"00110100011",
"00100101011",
"00111011111",
"00110100001",
"00111001010",
"00110001011",
"00111100001",
"00110011000",
"00100000110",
"00110110001",
"00110001110",
"00110010100",
"01000010100",
"00110001101",
"00101000001",
"00100101101",
"01000001110",
"00110111110",
"00110001011",
"00110011001",
"00101001001",
"00100100000",
"00111010110",

"00111000100",
"00110011000",
"00100011111",
"00101001011",
"00110100101",
"00110100001",
"00101001111",
"00101010101",
"00111000110",
"00010110100",
"00100001110",
"00101100001",
"00110011110",
"00110101101",
"00111100001",
"00100101110",
"00011010110",
"00110011100",
"00010010111",
"00100110011",
"00110110100",
"00110011011",
"00100101011",
"00101001000",
"00010110111",
"00100010001",
"00100011001",
"00010101011",
"00110100110",
"00101000111",
"00110010001",
"00101001010",
"01000101001",
"00011010110",
"00100101010",
"00010110101",
"00110001001",
"00110001010",
"00110111000",
"00110010101",
"00100011101",
"00101001100",
"00100111011",
"00110011010",
"00100111111",
"00100101111",
"00111001100",
"00100110110",
"00101011111",
"00110101010",
"00011011110",
"00011010011",
"00100101010",
"00110001010",
"00110100111",
"00110110101",
"00010110111",
"00101010101",
"00111011010",
"00110111111",
"00110101100",
"00110011101",
"00110000000",
"00101010010",
"00011100011",
"00110100111",
"00111011000",
"00100100111",
"00100110001",
"00100101000",
"00011100011",
"00100011011",
"00101001101",
"00101010101",
"00001011111",
"00011001000",
"00110110101",
"00110011100",
"00100010110",
"00110001100",
"00100111000",
"00101011110",
"00101000111",
"00111000101",
"00110000110",
"00011010101",
"00110001111",
"00101011101",
"00101000011",
"00110010101",
"00101001101",
"00100011001",
"00100101100",
"01000000010",
"00110111101",
"00100111100",
"00110011000",
"00100001110",
"00100010111",
"00111001101",

"00111000011",
"00101000110",
"00100011001",
"00100101111",
"00100111100",
"00101100000",
"00100110111",
"00101000111",
"00101010100",
"00010011101",
"00011000011",
"00100111100",
"00110001010",
"00100010111",
"00011000011",
"00100001101",
"00011010101",
"00101010111",
"00010010001",
"00011000000",
"00110101010",
"00110001010",
"00010010001",
"00100000110",
"00010110010",
"00100000011",
"00100010100",
"00010101001",
"00100110001",
"00100101010",
"00101011000",
"00100101111",
"00110001001",
"00010100010",
"00100001110",
"00010000101",
"00101000010",
"00101000000",
"00110100100",
"00110010011",
"00100011001",
"00010100110",
"00100101100",
"00101011001",
"00100000011",
"00011100010",
"00110011100",
"00011010111",
"00101011100",
"00100000110",
"00011001101",
"00010101011",
"00011100001",
"00110001000",
"00110100010",
"00100110001",
"00010110110",
"00100100011",
"00110100101",
"00110001011",
"00110011100",
"00101100011",
"00100110101",
"00100110111",
"00011010010",
"00101000010",
"00111000001",
"00011011011",
"00100101110",
"00010110000",
"00010011001",
"00100001101",
"00101001010",
"00101010100",
"00000111000",
"00010010010",
"00101010010",
"00101000100",
"00100010010",
"00110000010",
"00100110101",
"00100100001",
"00100111101",
"00100101010",
"00100111100",
"00010110101",
"00101100010",
"00100101100",
"00100011101",
"00110000110",
"00100011011",
"00100001100",
"00100011010",
"00100101010",
"00110110010",
"00100010111",
"00101000000",
"00011000000",
"00100010100",
"00110000111",

"00111000010",
"00100110100",
"00010110001",
"00100101101",
"00010000100",
"00100110111",
"00001011001",
"00100011010",
"00100100101",
"00010000011",
"00010001010",
"00010110010",
"00100000100",
"00010011011",
"00010101000",
"00010111101",
"00010001101",
"00100110000",
"00001000011",
"00010111010",
"00100110001",
"00100101011",
"00001010010",
"00010111010",
"00010011100",
"00001010101",
"00011000101",
"00001010010",
"00100101100",
"00011011111",
"00100111110",
"00100101001",
"00101011000",
"00010011001",
"00100000011",
"00000111000",
"00100001110",
"00100111101",
"00110011001",
"00110010001",
"00010001101",
"00010001100",
"00011011011",
"00101010000",
"00011011011",
"00010100001",
"00100111110",
"00010100100",
"00101000101",
"00011011110",
"00011000011",
"00010000110",
"00011010001",
"00101100001",
"00110010110",
"00100010001",
"00001100011",
"00100010101",
"00010111101",
"00101011100",
"00100110111",
"00011010101",
"00100100111",
"00100100001",
"00010101110",
"00100111110",
"00110010010",
"00010010111",
"00100100010",
"00010010111",
"00010001100",
"00010111011",
"00011000100",
"00010011101",
"00000110111",
"00010000110",
"00011000010",
"00100101010",
"00100000111",
"00010111101",
"00100100011",
"00010100111",
"00011010000",
"00100000000",
"00011100000",
"00010110100",
"00100001100",
"00010101100",
"00010101001",
"00101001011",
"00010000111",
"00100000010",
"00011001001",
"00100000001",
"00101100001",
"00011010110",
"00100101100",
"00010111010",
"00100000100",
"00011010001",

"00101100010",
"00100110010",
"00001011110",
"00011010101",
"00000111001",
"00100101000",
"00000101101",
"00011011101",
"00010010110",
"00001011110",
"00001011001",
"00010001000",
"00001100000",
"00001100010",
"00001001010",
"00010011110",
"00010000101",
"00011001010",
"00000110111",
"00010110111",
"00010100010",
"00100101001",
"00000011000",
"00010100110",
"00010010100",
"00001010001",
"00010100101",
"00001000100",
"00100001101",
"00010111101",
"00100011100",
"00100000110",
"00101001011",
"00001001100",
"00010111110",
"00000110010",
"00100000110",
"00100100111",
"00100011101",
"00100000111",
"00001010101",
"00001001001",
"00010001011",
"00100101110",
"00000011001",
"00010001010",
"00100111011",
"00010100011",
"00100101000",
"00010101110",
"00010111011",
"00000100010",
"00010011110",
"00100011000",
"00110001000",
"00011011101",
"00001000000",
"00010001011",
"00001011101",
"00100111001",
"00100000010",
"00011000001",
"00010110010",
"00100011100",
"00010100101",
"00001010110",
"00101011010",
"00010001001",
"00010111110",
"00010001101",
"00000111000",
"00010111010",
"00001011000",
"00001011110",
"00000100101",
"00001001110",
"00001011011",
"00100000011",
"00011010111",
"00010100111",
"00011001001",
"00010100000",
"00010001101",
"00010111011",
"00010111001",
"00010100011",
"00010110101",
"00010011010",
"00010000010",
"00100000111",
"00001100000",
"00010111100",
"00011000110",
"00011100011",
"00101010000",
"00010111000",
"00010100101",
"00010110011",
"00011010101",
"00010001001",

"00101011110",
"00010101100",
"00001001111",
"00010100010",
"00000101000",
"00011011001",
"00000100001",
"00001010000",
"00001001101",
"00000110000",
"00000100010",
"00000001000",
"00000111001",
"00000111011",
"00001000101",
"00001100000",
"00001011100",
"00010010000",
"00000010100",
"00001001001",
"00010100001",
"00000111010",
"00000010001",
"00000110111",
"00001100000",
"00000110111",
"00001010001",
"00000111111",
"00010111001",
"00010000011",
"00010110011",
"00011010101",
"00100101101",
"00000111100",
"00001010100",
"00000011110",
"00011011000",
"00010000000",
"00001000001",
"00000111100",
"00001010010",
"00001000101",
"00001000000",
"00011001100",
"00000010111",
"00000111100",
"00000100110",
"00010010100",
"00100001111",
"00010001111",
"00010100101",
"00000001100",
"00010001110",
"00000011000",
"00010100100",
"00011001011",
"00000110001",
"00000101001",
"00001001010",
"00100110111",
"00000110011",
"00010110101",
"00000011001",
"00010100101",
"00000010110",
"00000010101",
"00100011010",
"00000111100",
"00010101111",
"00000110111",
"00000010100",
"00000101011",
"00001010100",
"00001001110",
"00000011100",
"00000111000",
"00001010101",
"00010111100",
"00010100001",
"00010100011",
"00000111011",
"00000111101",
"00010000110",
"00000001001",
"00010010100",
"00001000111",
"00010101111",
"00010010100",
"00000111111",
"00010011100",
"00000011101",
"00000001010",
"00011000000",
"00010001110",
"00001011010",
"00010010110",
"00000110001",
"00010011101",
"00010010110",
"00001011010",

"00010100000",
"00000000100",
"00000011001",
"00000101100",
"00000001110",
"00011000110",
"00000011100",
"00000100001",
"00000111110",
"00000011001",
"00000011011",
"00000000001",
"00000011100",
"00000001001",
"00000100001",
"00000000101",
"00001011011",
"00000010010",
"00000001010",
"00001000100",
"00010000110",
"00000110000",
"00000000100",
"00000011010",
"00001011001",
"00000011101",
"00000010010",
"00000110001",
"00000110100",
"00000001111",
"00001000100",
"00010000010",
"00001001100",
"00000110100",
"00000100011",
"00000011101",
"00000000110",
"00001100010",
"00000100110",
"00000100011",
"00001001010",
"00000110101",
"00000101101",
"00010111101",
"00000000111",
"00000010010",
"00000011001",
"00010000011",
"00001000101",
"00010001110",
"00010011010",
"00000000100",
"00000001011",
"00000000110",
"00001011010",
"00010011110",
"00000001000",
"00000100110",
"00000101001",
"00011000101",
"00000100110",
"00000111001",
"00000000101",
"00010011000",
"00000001000",
"00000010100",
"00011011100",
"00000000111",
"00000011001",
"00000001011",
"00000001101",
"00000001101",
"00000111111",
"00000010011",
"00000011000",
"00000010111",
"00000111110",
"00000101001",
"00000001011",
"00000101010",
"00000011000",
"00000000101",
"00001001001",
"00000000000",
"00000110100",
"00000010101",
"00010101100",
"00010010010",
"00000000000",
"00001000101",
"00000000001",
"00000001000",
"00001010010",
"00000001000",
"00000011110",
"00000000011",
"00000101001",
"00001000011",
"00000011001",
"00000001001",


"10000111110",
"10000110001",
"10000110010",
"10000111010",
"10001001001",
"10000110101",
"10001000111",
"10000110111",
"10000100001",
"10001001110",
"10000110100",
"10001000101",
"10001001100",
"10000110101",
"10000100010",
"10000110000",
"10000001110",
"10001000100",
"10001001001",
"10001000010",
"10000100001",
"10000101011",
"10000111110",
"10000100011",
"10000010111",
"10000101010",
"10000111010",
"10001000011",
"10000011001",
"10000100100",
"10000111110",
"10000011001",
"10001010000",
"10000111011",
"10001001100",
"10000111011",
"10001000000",
"10000011100",
"10000010110",
"10001001110",
"10000011011",
"10000010011",
"10000111110",
"10001001110",
"10000100000",
"10000101101",
"10000101000",
"10000111110",
"10000010101",
"10001001111",
"10000110101",
"10001001111",
"10000111010",
"10000100111",
"10001000101",
"10001000111",
"10000111100",
"10001010010",
"10000111100",
"10001001000",
"10000110000",
"10001000110",
"10000101000",
"10000011101",
"10001001110",
"10000100110",
"10001010010",
"10001001000",
"10001000100",
"10000110110",
"10001010010",
"10000100111",
"10000010110",
"10001010000",
"10000100010",
"10001001101",
"10000011111",
"10000010011",
"10001000111",
"10000100100",
"10001000011",
"10000101011",
"10001001110",
"10001000100",
"10001000110",
"10001000101",
"10000110010",
"10000110000",
"10000111111",
"10001001111",
"10000111000",
"10000101100",
"10000111010",
"10001000101",
"10000110110",
"10000100010",
"10000110000",
"10000100100",
"10001001101",
"10001001010",

"10000100011",
"10000101110",
"10000001101",
"10000010010",
"10000111011",
"10000010110",
"10000100011",
"10000100100",
"10000010111",
"10001001010",
"10000001000",
"10000111110",
"10001000011",
"10000001111",
"10000011010",
"10000100111",
"10000001101",
"10001000001",
"10000011110",
"10000111000",
"10000011110",
"10000001100",
"10000010000",
"10000011010",
"10000001001",
"10000100111",
"10000100001",
"10000010100",
"10000001110",
"10000011111",
"10000110101",
"10000010011",
"10000111111",
"10000101100",
"10000001110",
"10000101001",
"10000110101",
"10000010100",
"10000001111",
"10000110111",
"10000010011",
"10000001111",
"10000100010",
"10000001101",
"10000010111",
"10000100010",
"10000100110",
"10000010111",
"10000000111",
"10001001110",
"10000010000",
"10001001110",
"10000001011",
"10000100101",
"10000001011",
"10000111010",
"10000000111",
"10001001101",
"10000001110",
"10000101000",
"10000100100",
"10000001100",
"10000001101",
"10000011010",
"10000101001",
"10000000101",
"10000010011",
"10000110110",
"10000110111",
"10000001001",
"10000110101",
"10000001000",
"10000000111",
"10001000011",
"10000011011",
"10001000010",
"10000010000",
"10000010000",
"10000001110",
"10000010110",
"10000101100",
"10000001000",
"10000111111",
"10000111100",
"10000010000",
"10000011101",
"10000100111",
"10000011000",
"10000100000",
"10000111010",
"10000100010",
"10000101011",
"10000010110",
"10000010000",
"10000010011",
"10000011110",
"10000010111",
"10000000111",
"10000101010",
"10000011001",

"01001011011",
"00110111110",
"01001100010",
"01000101011",
"01000010101",
"01000101101",
"01000010111",
"01001001101",
"01000101001",
"01001010110",
"01001011011",
"01000111001",
"01001010100",
"01000110010",
"01000001101",
"01000100000",
"01000001110",
"01000110100",
"01001100000",
"01001000111",
"01000100101",
"01001010010",
"01001011010",
"01001001101",
"01000110000",
"00111001111",
"01001011000",
"01001100001",
"01001011101",
"01001000010",
"01001100001",
"00100011101",
"01001001110",
"01000110111",
"01001011001",
"00110011001",
"01001001101",
"01000101110",
"01001010111",
"01001100011",
"01001001111",
"01000010010",
"01000010010",
"01000001011",
"01000100000",
"01001010001",
"01000111100",
"01001001101",
"00111000101",
"01001010000",
"01001010110",
"01001001001",
"01001010010",
"01001010000",
"01000110001",
"01000110111",
"01001001001",
"01000111101",
"01001011101",
"01001000000",
"01001000110",
"01001001000",
"01000000001",
"01001010101",
"01001001000",
"01000001111",
"01001000011",
"01001000010",
"01000111011",
"01000110101",
"01000101001",
"01001001100",
"01000101000",
"01000001000",
"01000010101",
"01000100000",
"01001011010",
"01000110000",
"01000011000",
"01000011111",
"01001000101",
"01000100000",
"01001010010",
"01000111011",
"01001100010",
"01001011101",
"01001011001",
"00110111100",
"01001010011",
"01000110110",
"01001010111",
"01000000010",
"01000110100",
"01001011011",
"01001011101",
"01000010111",
"01001010000",
"01000010110",
"01001011101",
"01001100011",

"01001010111",
"00110110011",
"00110010100",
"01000010011",
"00111011000",
"01000100011",
"00111100001",
"00111100000",
"01000010111",
"00110111101",
"01000010010",
"01000000101",
"01000011001",
"01000010011",
"00111000001",
"01000001000",
"01000001011",
"01000000011",
"01001011000",
"01001000100",
"00111000011",
"01000110111",
"01001010111",
"01000100100",
"01000010000",
"00111000111",
"01000011111",
"01000111001",
"01001010000",
"01000000110",
"01000100100",
"00011100010",
"01000100001",
"01000110100",
"01000110001",
"00110010011",
"01000001000",
"01000010100",
"01000110101",
"00111001101",
"01000101000",
"01000010000",
"00110011011",
"00101011001",
"00111011100",
"01000111101",
"01000100101",
"01000100011",
"00110111000",
"01000111001",
"01000001010",
"01000101001",
"00111000010",
"00111010001",
"01000001110",
"01000110010",
"01001000100",
"00110001000",
"01001010010",
"01000011001",
"01000111111",
"01000001101",
"00111010010",
"01000011001",
"01001000010",
"01000000111",
"00110110110",
"01000111000",
"00110011011",
"00011001000",
"00110110100",
"00111011110",
"01000010110",
"00110001101",
"01000001100",
"00110001000",
"01001010110",
"01000101000",
"01000010101",
"01000001011",
"00111000111",
"00110001000",
"01001001001",
"01000100110",
"01000010000",
"01000110000",
"01000100111",
"00100111101",
"01001001011",
"00110111011",
"01000110110",
"00111011000",
"01000100010",
"01001001010",
"01000111010",
"01000000100",
"01001001100",
"00110011100",
"01000010000",
"01000111110",

"00111011001",
"00110101100",
"00110000011",
"01000010010",
"00111001001",
"00110010110",
"00111001100",
"00110100001",
"00111011000",
"00110011000",
"00111000101",
"00111000000",
"01000010011",
"00111010111",
"00110101101",
"00110000111",
"00110100101",
"00110011100",
"01000100011",
"01000011001",
"00111000001",
"01000110100",
"01000100010",
"01000010001",
"01000001011",
"00110001011",
"00111001010",
"01000110001",
"01000010011",
"00110001001",
"01000000110",
"00011010010",
"01000010010",
"01000101111",
"01000001101",
"00101001000",
"00110000101",
"00111100001",
"00101001110",
"00110110101",
"01000100011",
"00101010101",
"00110001101",
"00101001011",
"00111001111",
"01000011000",
"01000011001",
"01000100001",
"00101010001",
"00110111010",
"00111001010",
"01000011000",
"00101011100",
"00101000110",
"00110011000",
"00111011100",
"01000101001",
"00101011001",
"01000011010",
"01000010100",
"01000000000",
"00111000000",
"00110111000",
"00111011000",
"00111001010",
"00111000101",
"00110000101",
"01000101110",
"00110001100",
"00010110011",
"00110110001",
"00110100000",
"00111001001",
"00101011011",
"00111011110",
"00101100011",
"01000111001",
"01000100011",
"00110100000",
"01000000010",
"00111000110",
"00110000110",
"01000000000",
"00101010100",
"00111011000",
"00011000110",
"01000001110",
"00100110100",
"00110100100",
"00101010000",
"00111010001",
"00110101010",
"01000011010",
"01000000000",
"01000010001",
"00110110100",
"01000100101",
"00101011111",
"00101000011",
"00101000100",

"00111010101",
"00100001100",
"00101011011",
"01000000001",
"00110101010",
"00110001001",
"00101010111",
"00110001001",
"00110110011",
"00100111011",
"00110101111",
"00110101010",
"00110110111",
"00101000010",
"00110101100",
"00101000110",
"00110011101",
"00100111101",
"00111011000",
"00111011110",
"00110110000",
"00111010011",
"00110000110",
"00111010011",
"00111100010",
"00110000011",
"00100011010",
"01000110000",
"00111011011",
"00110000001",
"00101010111",
"00010101001",
"00101010101",
"00101000111",
"00111100010",
"00100001101",
"00110000001",
"00101100000",
"00100000001",
"00110100101",
"01000011011",
"00100011101",
"00110001000",
"00101000110",
"00110110000",
"00111010011",
"00111011011",
"01000001110",
"00100110111",
"00110110110",
"00101011100",
"00110100111",
"00100110100",
"00101000011",
"00100111111",
"00111001100",
"00101011001",
"00100010100",
"00111100010",
"00101100001",
"00101011110",
"00110000010",
"00110100001",
"00111010010",
"00111000100",
"00110100100",
"00110000011",
"00110101100",
"00101010011",
"00010101010",
"00110010000",
"00101011111",
"00110101111",
"00100001101",
"00110101111",
"00100100000",
"01000011011",
"00100010100",
"00110001010",
"00111000110",
"00110110010",
"00101010100",
"00101011100",
"00100110011",
"00110001011",
"00011000101",
"00111010001",
"00100110000",
"00101100000",
"00011100010",
"00110101100",
"00110011110",
"00110011100",
"00111010100",
"00111100001",
"00110000000",
"01000000001",
"00101000100",
"00100110110",
"00100110110",

"00111001110",
"00011100001",
"00101010001",
"00110101101",
"00110011110",
"00100011011",
"00101000101",
"00101011101",
"00101010101",
"00011010100",
"00110010100",
"00110010000",
"00110100110",
"00100010100",
"00010100110",
"00100010101",
"00011011110",
"00100101111",
"00110111110",
"00100101011",
"00100010001",
"00110011101",
"00100101011",
"00110111111",
"00101100011",
"00101000001",
"00100010100",
"00111010110",
"00110011110",
"00101000001",
"00010101111",
"00010011111",
"00101010010",
"00100011000",
"00101000110",
"00011100001",
"00100011100",
"00100101111",
"00010100110",
"00110011000",
"00100100101",
"00100011100",
"00100111001",
"00101000011",
"00101100010",
"00110110100",
"00111001100",
"00110000010",
"00100010101",
"00110100110",
"00101011000",
"00110001010",
"00100010101",
"00100000011",
"00011010011",
"00100001011",
"00011001011",
"00011011011",
"00111100000",
"00100011110",
"00101000011",
"00101000111",
"00101010111",
"00100110111",
"00110101011",
"00101001110",
"00110000001",
"00110000111",
"00001011001",
"00010001001",
"00011011100",
"00101001111",
"00110001100",
"00010110001",
"00110011100",
"00100010001",
"00111000101",
"00011100001",
"00011010111",
"00110010100",
"00110010101",
"00011011101",
"00100001101",
"00100110010",
"00110000001",
"00010110010",
"00100101100",
"00100101000",
"00100011110",
"00010110100",
"00110000011",
"00110011101",
"00101011010",
"00110111111",
"00111010011",
"00100101001",
"00110111111",
"00100111010",
"00010011000",
"00100011111",

"00110100101",
"00011001010",
"00101000000",
"00100001010",
"00110011100",
"00010101011",
"00100100101",
"00101010001",
"00100110011",
"00010110111",
"00110000100",
"00101001101",
"00110001100",
"00010111011",
"00010011000",
"00010001100",
"00010100001",
"00010010101",
"00110111100",
"00011011110",
"00010100111",
"00100011101",
"00001011011",
"00101001100",
"00101100010",
"00100110010",
"00100000110",
"00110111011",
"00110000011",
"00100111101",
"00010001100",
"00010011010",
"00101000011",
"00011010000",
"00100110100",
"00011010011",
"00100010001",
"00011010100",
"00001010110",
"00100110001",
"00011011001",
"00011001001",
"00100100010",
"00101000010",
"00100011111",
"00100110000",
"00100011010",
"00011000010",
"00100001000",
"00110011011",
"00100001000",
"00101000101",
"00011011001",
"00011000101",
"00010101110",
"00100000110",
"00010101011",
"00011001110",
"00111011100",
"00100011010",
"00100010011",
"00011011010",
"00011011110",
"00100001111",
"00110010010",
"00101000001",
"00101100011",
"00101100010",
"00001001111",
"00001011010",
"00010011011",
"00101000110",
"00110001001",
"00010100000",
"00101001001",
"00011011000",
"00110100010",
"00011001000",
"00010000011",
"00110000111",
"00110001001",
"00010110011",
"00011001001",
"00100011100",
"00100110101",
"00010101010",
"00010011111",
"00011011100",
"00010101101",
"00010110001",
"00100001110",
"00010101111",
"00010110011",
"00110100001",
"00111000100",
"00100001100",
"00100110101",
"00100101101",
"00010010011",
"00100011100",

"00100110000",
"00010001001",
"00100000111",
"00011001010",
"00101010000",
"00010010010",
"00010001010",
"00010001100",
"00100101101",
"00010011010",
"00100001110",
"00100001101",
"00110000100",
"00010000001",
"00001011010",
"00010000100",
"00010001110",
"00010010000",
"00100010010",
"00011011000",
"00010000011",
"00010011101",
"00001001011",
"00100111111",
"00010101010",
"00100100011",
"00011011111",
"00110011101",
"00100011010",
"00011000011",
"00001100000",
"00010000101",
"00100100001",
"00010111110",
"00100000111",
"00010010000",
"00100001110",
"00010100001",
"00000110110",
"00100010000",
"00011010010",
"00011000110",
"00100001110",
"00100110110",
"00011100000",
"00011001011",
"00100000100",
"00010101000",
"00100000110",
"00110011000",
"00010101010",
"00100100100",
"00001011111",
"00000101001",
"00010001000",
"00010110110",
"00010001100",
"00010110001",
"00011000111",
"00010111100",
"00011011010",
"00011001000",
"00011010111",
"00011001101",
"00110001111",
"00100101100",
"00101011011",
"00101001000",
"00001001110",
"00001010110",
"00001000111",
"00010110111",
"00100110001",
"00001100011",
"00100101011",
"00011010101",
"00101000101",
"00010010110",
"00001011010",
"00100011011",
"00101010111",
"00010110010",
"00001010010",
"00011011000",
"00100001110",
"00010000101",
"00010000010",
"00011001110",
"00010010001",
"00001011101",
"00011000010",
"00010011011",
"00010011011",
"00110001110",
"00011010010",
"00011001111",
"00011011001",
"00100011010",
"00000011110",
"00011001011",

"00011000001",
"00001010000",
"00010111101",
"00011000001",
"00101000001",
"00010001000",
"00001100010",
"00010001011",
"00100010011",
"00010000000",
"00010011100",
"00000111000",
"00011000011",
"00001100001",
"00001001011",
"00001011111",
"00001010100",
"00010000010",
"00011010100",
"00010111111",
"00001010001",
"00010000011",
"00000110001",
"00010111111",
"00001011001",
"00011010001",
"00000111110",
"00100111010",
"00011100011",
"00010111011",
"00001010110",
"00010000001",
"00010001101",
"00001100011",
"00011010010",
"00010000110",
"00100000100",
"00010011010",
"00000101110",
"00011010010",
"00010001010",
"00001010100",
"00001000110",
"00100100000",
"00011011010",
"00010011010",
"00010111010",
"00010001000",
"00010101011",
"00100001100",
"00001001110",
"00010100000",
"00001010100",
"00000011111",
"00000100010",
"00010011000",
"00010001011",
"00010000000",
"00001010101",
"00001011110",
"00010111010",
"00010000100",
"00001001011",
"00001011011",
"00101000010",
"00010100100",
"00101010001",
"00010011111",
"00000011010",
"00000111001",
"00000101110",
"00010101111",
"00100100111",
"00000111001",
"00010110111",
"00010100110",
"00100100010",
"00010010001",
"00000010010",
"00100001100",
"00100011001",
"00001010010",
"00001000110",
"00010111001",
"00011000010",
"00001010111",
"00001100000",
"00010101110",
"00010000001",
"00001000010",
"00010010100",
"00001011010",
"00010000001",
"00100111011",
"00001100010",
"00010101111",
"00011010100",
"00010100011",
"00000011011",
"00010100101",

"00000100101",
"00000010001",
"00010000100",
"00010101100",
"00100111101",
"00000100100",
"00000110100",
"00000110001",
"00010100000",
"00000101110",
"00001000100",
"00000101110",
"00001011111",
"00000011100",
"00000111010",
"00000110000",
"00001000100",
"00000100110",
"00010010000",
"00001010010",
"00001001001",
"00000010011",
"00000100110",
"00001011101",
"00001001100",
"00010100111",
"00000101011",
"00010011000",
"00011000000",
"00010110000",
"00000011001",
"00000101110",
"00001010111",
"00001001001",
"00010101100",
"00000111011",
"00011001010",
"00001010001",
"00000101011",
"00010000110",
"00001010011",
"00001001000",
"00000010100",
"00100000100",
"00010101010",
"00001011110",
"00010011100",
"00000100100",
"00000101011",
"00001010101",
"00000010000",
"00000111111",
"00001001000",
"00000011101",
"00000011010",
"00001001011",
"00001100000",
"00000101011",
"00000011111",
"00000110001",
"00001011000",
"00001000010",
"00000111111",
"00001001001",
"00010011010",
"00001001001",
"00011011001",
"00010000010",
"00000010110",
"00000110010",
"00000101010",
"00010000010",
"00100010100",
"00000101101",
"00010101010",
"00001011001",
"00100000110",
"00000011001",
"00000000100",
"00100000010",
"00011010100",
"00000111111",
"00000110100",
"00000111000",
"00010011111",
"00000110000",
"00001010100",
"00010100100",
"00000110000",
"00000001110",
"00001001011",
"00001010000",
"00000100010",
"00100011110",
"00000011001",
"00010011010",
"00011001001",
"00010010000",
"00000010011",
"00010011000",

"00000011111",
"00000000001",
"00001100010",
"00000010111",
"00100001111",
"00000000010",
"00000101000",
"00000100001",
"00010000011",
"00000010001",
"00000000011",
"00000011010",
"00000110011",
"00000000001",
"00000100010",
"00000100110",
"00000000100",
"00000000010",
"00000011000",
"00000010001",
"00000010000",
"00000010010",
"00000100011",
"00000111010",
"00000111100",
"00000101111",
"00000010110",
"00000001010",
"00010011000",
"00010010001",
"00000001101",
"00000000010",
"00000011111",
"00000110100",
"00000101001",
"00000001011",
"00011000100",
"00000100000",
"00000011110",
"00000100001",
"00000010011",
"00000111111",
"00000000101",
"00010011000",
"00001011101",
"00000001001",
"00010001111",
"00000001011",
"00000010010",
"00000000010",
"00000000101",
"00000010100",
"00001000110",
"00000000011",
"00000001000",
"00000110101",
"00000011011",
"00000001111",
"00000010111",
"00000100110",
"00000011111",
"00000100100",
"00000010001",
"00001000001",
"00000100000",
"00000010001",
"00010001111",
"00000000111",
"00000000101",
"00000001111",
"00000001111",
"00010000000",
"00010110001",
"00000000000",
"00000000101",
"00000111101",
"00010011110",
"00000010111",
"00000000001",
"00000100101",
"00010111001",
"00000001101",
"00000000010",
"00000100111",
"00010001100",
"00000010011",
"00000000000",
"00000001010",
"00000001000",
"00000000101",
"00000110101",
"00001001110",
"00000000100",
"00000110111",
"00000010001",
"00010000101",
"00011000001",
"00000000101",
"00000001110",
"00010010000",


"10000110111",
"10001000000",
"10001000000",
"10001000100",
"10000110001",
"10001000010",
"10000101101",
"10000111101",
"10000010001",
"10001000111",
"10001000001",
"10000101010",
"10000110101",
"10001010001",
"10001001011",
"10000111111",
"10001001111",
"10000101000",
"10000100010",
"10001000011",
"10001000010",
"10001000011",
"10001001110",
"10000101011",
"10000110010",
"10001001000",
"10001010001",
"10001010000",
"10001000010",
"10000101010",
"10001001010",
"10001000001",
"10000111101",
"10001010010",
"10000101110",
"10001001010",
"10001001100",
"10000100010",
"10001000111",
"10001000100",
"10001000000",
"10000111010",
"10001001011",
"10000101100",
"10001000010",
"10000011001",
"10000111000",
"10001000111",
"10001001100",
"10001010001",
"10001000011",
"10001001111",
"10000111111",
"10001001010",
"10000100101",
"10001000101",
"10001001100",
"10000101011",
"10001001100",
"10000110010",
"10001001011",
"10000101001",
"10000101110",
"10001000001",
"10000111011",
"10001001111",
"10000110100",
"10000100111",
"10001010001",
"10001000000",
"10001001010",
"10000011110",
"10000110101",
"10001001100",
"10000101001",
"10001000111",
"10000100101",
"10001000011",
"10001000001",
"10000010111",
"10001001111",
"10000110110",
"10000111110",
"10000100011",
"10000111101",
"10000110001",
"10000100100",
"10000110110",
"10000111001",
"10000111001",
"10001000111",
"10000011101",
"10001001011",
"10000110011",
"10000101111",
"10000110101",
"10001000111",
"10000100100",
"10000011110",
"10001001000",

"10000110000",
"10000111000",
"10000011110",
"10000010110",
"10000011000",
"10000111010",
"10000010100",
"10000010010",
"10000001100",
"10000111101",
"10000010010",
"10000001010",
"10000100000",
"10000110010",
"10001001010",
"10000011100",
"10000010110",
"10000010001",
"10000011000",
"10000001111",
"10000101011",
"10000010001",
"10000111010",
"10000100111",
"10000001010",
"10000110110",
"10000001101",
"10000011011",
"10000000110",
"10000010000",
"10000001011",
"10000101100",
"10000011110",
"10000010010",
"10000010111",
"10000100011",
"10000110000",
"10000010100",
"10000011110",
"10000111000",
"10000110001",
"10000101000",
"10000100010",
"10000100100",
"10000100111",
"10000010101",
"10000000101",
"10000001111",
"10001000010",
"10000000110",
"10000001101",
"10000110011",
"10000110000",
"10000101101",
"10000010110",
"10000001111",
"10000110111",
"10000001101",
"10000011001",
"10000011101",
"10001000110",
"10000010110",
"10000100100",
"10000100111",
"10000011011",
"10000011111",
"10000110011",
"10000010001",
"10001010000",
"10000111000",
"10000101011",
"10000011101",
"10000100100",
"10000110101",
"10000011001",
"10000110110",
"10000011101",
"10000001110",
"10000010100",
"10000001011",
"10000011010",
"10000010110",
"10000101001",
"10000011101",
"10000001011",
"10000100110",
"10000100000",
"10000101111",
"10000001000",
"10000010001",
"10000001101",
"10000010010",
"10001001000",
"10000001010",
"10000010000",
"10000010011",
"10000001111",
"10000001010",
"10000010000",
"10001000011",

"01001000000",
"01001011101",
"01001000011",
"01000110010",
"01000100001",
"01001010011",
"01000010001",
"01000101100",
"01001100010",
"01000100011",
"01000001011",
"01001010101",
"01000001100",
"01000011110",
"01001000011",
"01000110001",
"01001000101",
"00111011111",
"01001001000",
"01000111110",
"01001100000",
"01001010011",
"01001010100",
"01001000111",
"01000111001",
"01001100010",
"01001011010",
"01000001100",
"01001100010",
"01000011011",
"01001011010",
"01001010011",
"01001100001",
"01001010001",
"01001001111",
"01001011001",
"01000111101",
"01000000101",
"01001011011",
"00111001111",
"00110011110",
"01001010000",
"01001000101",
"01001010111",
"01001100000",
"01000110000",
"01001010011",
"01001010110",
"01001011100",
"01001100011",
"01001011010",
"01000111011",
"01000110110",
"00111010011",
"01001000101",
"01001100011",
"01000101100",
"01000110001",
"01001010110",
"00111010101",
"01000111010",
"01000110011",
"01001100000",
"01000101101",
"01000111101",
"01000111111",
"01001000110",
"00111011011",
"01000101011",
"01000010011",
"01001001011",
"01001000100",
"01001011111",
"01000110000",
"01000110011",
"01000101111",
"01000010100",
"01001001001",
"01000110000",
"01001001010",
"01001010101",
"01001000101",
"00111010100",
"01001011100",
"01001010110",
"00111001011",
"01001010110",
"01000100011",
"01001100011",
"01001011111",
"01001011110",
"01000010111",
"01001011110",
"01000101101",
"01000101101",
"01001000011",
"01001000111",
"01001011000",
"01001000111",
"01000111101",

"01000111111",
"01001001101",
"01000111101",
"01000001110",
"01000010001",
"00110001100",
"00111010001",
"00111000010",
"01000101010",
"00111011000",
"01000000010",
"01001000010",
"00110111101",
"01000010100",
"01000110111",
"01000000110",
"01000101011",
"00111011000",
"01000010101",
"01000000101",
"01001010010",
"01000010111",
"01000111010",
"01000010011",
"01000010101",
"00101011011",
"01000111111",
"00111001000",
"01001010001",
"01000000001",
"00110100110",
"01000100011",
"00111001001",
"01000111011",
"01000000110",
"00111000000",
"01000011001",
"00111001100",
"01000110100",
"00110011100",
"00110000011",
"01000011110",
"01000111001",
"01000111010",
"01000110010",
"01000100110",
"01000000100",
"01000010010",
"01001010010",
"00110100011",
"01000101111",
"01000010100",
"01000011011",
"00111001000",
"01000111010",
"01001010100",
"01000100010",
"01000010110",
"01001001101",
"00111001010",
"01000111000",
"00110110000",
"01001001111",
"00111000100",
"00101001100",
"01000101010",
"01000011101",
"00110010010",
"00111001011",
"00111001000",
"01000101111",
"01001000011",
"01001011010",
"01000100111",
"01000101111",
"00111000110",
"00111100000",
"01001000111",
"01000001001",
"01000110110",
"01000110010",
"00111100001",
"00110001100",
"01000010110",
"01001000111",
"00110111100",
"01001010101",
"00101010111",
"01000000001",
"01001000100",
"01000110011",
"01000010110",
"01000101111",
"00110001111",
"00111011111",
"01000101111",
"01000101101",
"00111100000",
"01000111111",
"01000100011",

"01000001010",
"00110010010",
"00110011000",
"00110101011",
"00110111111",
"00101100010",
"00110110011",
"00110100001",
"00110100100",
"00110010001",
"00111011110",
"01000011101",
"00110110000",
"00101000110",
"00110011001",
"00111011001",
"00111010101",
"00110010001",
"00110111101",
"00111011011",
"01000110100",
"00111100011",
"01000110011",
"01000010010",
"01000010011",
"00101001100",
"00110001000",
"00101011001",
"01000101000",
"00111100001",
"00100111101",
"01000010110",
"00110001001",
"01000101001",
"00110101000",
"00110011000",
"01000010101",
"00110011110",
"00111010011",
"00101010101",
"00100000011",
"01000010100",
"00110111110",
"01000101111",
"00110101011",
"00111000100",
"00110111001",
"00110111001",
"00110010000",
"00110010111",
"01000000001",
"00111010110",
"01000010001",
"00111000001",
"00100101000",
"01000110011",
"01000001101",
"01000000000",
"00111100010",
"00110100101",
"01000110110",
"00110101100",
"01000110100",
"00111000001",
"00101000000",
"01000100011",
"00110011111",
"00110001010",
"00110011011",
"00111000110",
"01000100001",
"00110101101",
"00110111011",
"00110101000",
"00111001111",
"00110100000",
"00110010100",
"01000001000",
"01000000000",
"00111011111",
"00111011011",
"00111001111",
"00100100111",
"01000001001",
"00110110101",
"00110000111",
"01001000010",
"00100111011",
"00110110111",
"00110100111",
"01000100000",
"01000000000",
"01000100011",
"00100001011",
"00110001110",
"00111010001",
"01000101100",
"00110110111",
"01000111001",
"00111010001",

"00111011111",
"00110000001",
"00110010010",
"00110011010",
"00101000101",
"00101010100",
"00110101100",
"00110001010",
"00101001101",
"00110000111",
"00110011011",
"00111100011",
"00100110110",
"00100101001",
"00101011010",
"00100101101",
"00110101011",
"00100011110",
"00110001101",
"00110101011",
"01000011001",
"00110111111",
"01000100010",
"01000000110",
"01000001111",
"00100011010",
"00101011000",
"00100001111",
"00111000011",
"00100100110",
"00100110001",
"00110110101",
"00110000101",
"00101001111",
"00100101110",
"00101010110",
"00110110000",
"00110011000",
"00110101001",
"00101001011",
"00010001101",
"01000000110",
"00110101101",
"00111011010",
"00110100100",
"00110011000",
"00110110111",
"00101001010",
"00110001101",
"00110010110",
"00101011001",
"00101010000",
"00110010101",
"00110101110",
"00100010110",
"01000011100",
"00111001011",
"00110101111",
"00111010010",
"00110000111",
"01000011000",
"00100111010",
"01000001001",
"00110000110",
"00100111001",
"01000011010",
"00110011100",
"00010110111",
"00101100000",
"00110011010",
"01000001010",
"00110100000",
"00101000100",
"00110100010",
"00110110011",
"00101010100",
"00110010000",
"00110101000",
"00111100001",
"00110001111",
"00110011110",
"00110001100",
"00100000001",
"01000001000",
"00110101001",
"00110000010",
"01000011010",
"00011010101",
"00110011011",
"00110010111",
"01000000011",
"00100010100",
"01000001101",
"00100000110",
"00110001101",
"00111001000",
"01000001000",
"00110001010",
"01000011011",
"00110101011",

"00111010110",
"00101001100",
"00100100101",
"00100110001",
"00100100010",
"00100101110",
"00100100100",
"00110000000",
"00100000011",
"00100101010",
"00100010010",
"00111011010",
"00100110010",
"00100101000",
"00011010010",
"00100101010",
"00100001101",
"00100001000",
"00110001010",
"00110100101",
"00111100000",
"00110111000",
"01000011110",
"01000000010",
"00110101111",
"00010110100",
"00100100001",
"00011011000",
"00101010111",
"00100100101",
"00100100110",
"00101010111",
"00101011000",
"00100111000",
"00100101100",
"00101001101",
"00110101000",
"00101001000",
"00110100101",
"00011001110",
"00010001011",
"00111100001",
"00110010000",
"00110000011",
"00110100011",
"00101100010",
"00110110100",
"00100110101",
"00100111001",
"00110001101",
"00100011011",
"00101000111",
"00101010101",
"00110101011",
"00011100011",
"00101011001",
"00110010101",
"00011001011",
"00101011001",
"00101010110",
"01000010110",
"00100111000",
"00111010010",
"00101001111",
"00010110111",
"00110110111",
"00101011110",
"00010101011",
"00101011011",
"00101100011",
"00111100011",
"00110001001",
"00100101110",
"00101000101",
"00100111111",
"00100100111",
"00101011111",
"00101001100",
"00110000011",
"00110001100",
"00110001010",
"00101010100",
"00011001110",
"00111011001",
"00101011011",
"00101010001",
"00111010110",
"00011010100",
"00110001100",
"00010101011",
"00111011111",
"00100010000",
"01000000101",
"00011010110",
"00101100011",
"00111000000",
"01000000111",
"00100001111",
"01000001111",
"00110100010",

"00101001010",
"00010111001",
"00100100010",
"00100100010",
"00010000100",
"00100100101",
"00011001010",
"00101011001",
"00100000010",
"00011010100",
"00011001001",
"00110110110",
"00100100111",
"00100100101",
"00010101001",
"00010110011",
"00011000111",
"00010110110",
"00101000111",
"00101100010",
"00111000000",
"00100100100",
"01000010001",
"00111011111",
"00100001100",
"00010001011",
"00100010111",
"00010110101",
"00100101111",
"00100100100",
"00001011101",
"00100110001",
"00101010010",
"00100101100",
"00100001110",
"00101000001",
"00110100111",
"00001010000",
"00110011001",
"00011001101",
"00001011110",
"00110011011",
"00101100010",
"00101011001",
"00101001111",
"00100000101",
"00110001100",
"00011010110",
"00011011001",
"00100111111",
"00011011100",
"00011011010",
"00101010001",
"00110010010",
"00011010011",
"00101000100",
"00100010101",
"00010111011",
"00011001111",
"00101010100",
"00110100001",
"00011010101",
"00110111000",
"00100001100",
"00010100111",
"00110100011",
"00100110110",
"00010101010",
"00101001001",
"00011011111",
"00101100011",
"00100100000",
"00100011101",
"00100111110",
"00100111101",
"00100010101",
"00101001011",
"00100111011",
"00101001010",
"00100110000",
"00101000011",
"00101010010",
"00010100001",
"00110101111",
"00100010001",
"00100101011",
"00111010010",
"00011001101",
"00100010010",
"00000100001",
"00110101100",
"00011011110",
"00111100000",
"00011001011",
"00100110100",
"00110011111",
"00110011010",
"00100000111",
"00110111010",
"00110001110",

"00011011011",
"00001011101",
"00011010000",
"00011100011",
"00001010010",
"00010010001",
"00001000011",
"00100011000",
"00011000001",
"00010000001",
"00010001000",
"00110101101",
"00100010100",
"00010101000",
"00010000000",
"00010000110",
"00010001011",
"00010001000",
"00010010110",
"00100011111",
"00110011000",
"00010100010",
"01000001101",
"00110001011",
"00010010010",
"00001011110",
"00100010011",
"00001001111",
"00011010100",
"00011001000",
"00001001000",
"00011010011",
"00100110010",
"00010101101",
"00100001101",
"00100001011",
"00100000010",
"00001000111",
"00110010001",
"00010111101",
"00000100110",
"00100100011",
"00100111000",
"00100000010",
"00100100000",
"00011010100",
"00101010011",
"00011001001",
"00010111101",
"00010010010",
"00011000011",
"00011010111",
"00101000111",
"00101010110",
"00010111011",
"00011010101",
"00100000111",
"00001010011",
"00011001001",
"00100001010",
"00100101000",
"00010111011",
"00110011001",
"00100000100",
"00010100101",
"00101010111",
"00100001101",
"00010001000",
"00100101011",
"00010101011",
"00011000011",
"00011100011",
"00100001011",
"00100101101",
"00100001000",
"00010100001",
"00011011001",
"00100101110",
"00100101110",
"00100101100",
"00011011101",
"00100111000",
"00010001110",
"00010101100",
"00010100011",
"00011011111",
"00110000010",
"00010111001",
"00100001000",
"00000010100",
"00011001110",
"00011001000",
"00100000111",
"00011000100",
"00100101011",
"00101011011",
"00110011001",
"00100000101",
"00011010001",
"00100100110",

"00010101111",
"00000101011",
"00010101110",
"00010011111",
"00001001111",
"00000110010",
"00001000001",
"00011011000",
"00010100110",
"00010000000",
"00000110101",
"00110010100",
"00001001000",
"00010001011",
"00001011010",
"00001000111",
"00000110100",
"00001011001",
"00001011101",
"00011011111",
"00101010110",
"00010011010",
"01000000100",
"00011011000",
"00000101001",
"00000100000",
"00010010011",
"00000110110",
"00011000111",
"00010001100",
"00000100101",
"00010001011",
"00100000011",
"00010010100",
"00011000111",
"00011010100",
"00001001000",
"00000101011",
"00101001110",
"00010010100",
"00000100011",
"00011001111",
"00001001000",
"00011000011",
"00010001101",
"00010110111",
"00100001010",
"00010111011",
"00010101111",
"00010000011",
"00001010110",
"00000110001",
"00011011100",
"00101000010",
"00010101111",
"00001100001",
"00100000001",
"00001010001",
"00010010000",
"00011010111",
"00011011111",
"00001010111",
"00100101010",
"00011000111",
"00010011100",
"00101001110",
"00000110101",
"00010000001",
"00011000000",
"00001010110",
"00010101100",
"00011010010",
"00010110010",
"00011010111",
"00001001000",
"00001011011",
"00011001010",
"00010011001",
"00011010111",
"00010011001",
"00011010100",
"00100001101",
"00010001001",
"00010100100",
"00010011101",
"00010110011",
"00100101101",
"00001011100",
"00010100100",
"00000010001",
"00010100011",
"00011000110",
"00011011000",
"00001010100",
"00100010111",
"00100110101",
"00100011110",
"00011000110",
"00010110111",
"00011010011",

"00010001110",
"00000010000",
"00001001010",
"00001001011",
"00000100111",
"00000010001",
"00000111101",
"00000000110",
"00000111000",
"00000110000",
"00000101110",
"00100111011",
"00000001010",
"00001100011",
"00000101100",
"00001000000",
"00000101101",
"00001011000",
"00001001101",
"00010010100",
"00010010011",
"00010001000",
"00110001011",
"00010011111",
"00000011000",
"00000010100",
"00010001110",
"00000011100",
"00010011101",
"00000100001",
"00000100001",
"00001001111",
"00000111110",
"00010001011",
"00010001110",
"00010100111",
"00000111000",
"00000011100",
"00000110001",
"00001011010",
"00000010011",
"00010100000",
"00001000000",
"00010011100",
"00000111100",
"00001001110",
"00010100100",
"00010011000",
"00010001001",
"00000101100",
"00000111100",
"00000001010",
"00001001111",
"00100000100",
"00010010110",
"00001010000",
"00011011011",
"00000100101",
"00000101110",
"00010010101",
"00010101000",
"00000010110",
"00010100101",
"00011000100",
"00010000111",
"00000100000",
"00000011001",
"00001001001",
"00001011010",
"00001000111",
"00001100000",
"00010110110",
"00000111011",
"00010010101",
"00001000001",
"00001010110",
"00011000110",
"00010001000",
"00001100000",
"00001010111",
"00010110101",
"00001011010",
"00001100010",
"00010001010",
"00000010011",
"00001010001",
"00100100011",
"00000110111",
"00000110000",
"00000001110",
"00001010010",
"00000100010",
"00010101010",
"00001000001",
"00011001110",
"00010000111",
"00011010011",
"00010110000",
"00001001001",
"00010000010",

"00001100010",
"00000000001",
"00001000010",
"00000000001",
"00000000010",
"00000000101",
"00000100100",
"00000000011",
"00000010010",
"00000101111",
"00000010001",
"00100010100",
"00000001000",
"00001001011",
"00000101001",
"00000000100",
"00000100101",
"00000011000",
"00000000110",
"00001001011",
"00010001001",
"00000001010",
"00110001001",
"00000111011",
"00000000011",
"00000010001",
"00000001111",
"00000000010",
"00001001010",
"00000000010",
"00000010100",
"00000100011",
"00000011100",
"00001000100",
"00000110110",
"00000001100",
"00000000010",
"00000010011",
"00000000010",
"00000011000",
"00000010010",
"00010010111",
"00000000011",
"00000101111",
"00000000011",
"00000110010",
"00000001100",
"00000010100",
"00000110101",
"00000101011",
"00000011010",
"00000001001",
"00000000101",
"00000100001",
"00000100001",
"00001001010",
"00010011001",
"00000010001",
"00000101101",
"00000110110",
"00010000101",
"00000010010",
"00000110101",
"00010101000",
"00000011100",
"00000000011",
"00000000010",
"00000111111",
"00000101000",
"00000110011",
"00000010011",
"00010010100",
"00000110011",
"00000100001",
"00000111110",
"00000001001",
"00000001011",
"00001001101",
"00000100111",
"00001000000",
"00000101010",
"00000101111",
"00000101000",
"00000110100",
"00000001001",
"00000111001",
"00010101100",
"00000110100",
"00000010000",
"00000001100",
"00000100000",
"00000010011",
"00000101100",
"00000010011",
"00000100111",
"00000000101",
"00000110110",
"00001011000",
"00000011111",
"00000001001",


"10000110000",
"10000101001",
"10001001100",
"10001001000",
"10000101010",
"10000111000",
"10000111011",
"10001001011",
"10000111001",
"10000011101",
"10000111011",
"10001000111",
"10000110110",
"10000011001",
"10000011000",
"10001010001",
"10000011110",
"10001000100",
"10000111110",
"10000010101",
"10001001110",
"10001001101",
"10000110010",
"10000110001",
"10000011010",
"10000110011",
"10000110101",
"10001001001",
"10001000001",
"10001010000",
"10000111110",
"10001010000",
"10001001010",
"10001001010",
"10001000010",
"10000111000",
"10000011110",
"10001000111",
"10001000011",
"10000111100",
"10000110000",
"10000100111",
"10001001001",
"10001001100",
"10001001100",
"10001001101",
"10000011011",
"10000100110",
"10000111111",
"10000010101",
"10001010001",
"10000010111",
"10000111100",
"10001001001",
"10001000010",
"10001001001",
"10000110101",
"10001001000",
"10001010001",
"10000111110",
"10001010000",
"10000111110",
"10001001100",
"10000101110",
"10000111111",
"10001001101",
"10000100010",
"10000011110",
"10000011000",
"10000110001",
"10000111001",
"10000111011",
"10001001010",
"10000111011",
"10001000101",
"10000110011",
"10001001000",
"10001001101",
"10000111001",
"10000111000",
"10000011010",
"10000111011",
"10000111011",
"10001010010",
"10001001100",
"10001010010",
"10000011011",
"10001000001",
"10000011100",
"10000010010",
"10000110100",
"10001000101",
"10001001011",
"10000011011",
"10000101111",
"10001010010",
"10001001010",
"10001000100",
"10000111000",
"10000110100",

"10000100000",
"10000100110",
"10000001100",
"10000001111",
"10000011111",
"10000011010",
"10000001110",
"10000100001",
"10000110011",
"10000001111",
"10000101010",
"10001000110",
"10000100011",
"10000001010",
"10000010100",
"10001010000",
"10000010110",
"10000001000",
"10000011000",
"10000001110",
"10000010100",
"10000011000",
"10000011011",
"10000000111",
"10000011000",
"10000010101",
"10000010011",
"10000001100",
"10000001111",
"10001001101",
"10000001111",
"10000011101",
"10000011101",
"10000101010",
"10000010100",
"10000100101",
"10000010100",
"10001000110",
"10000000101",
"10000011110",
"10000100000",
"10000010010",
"10000001011",
"10000011000",
"10000101110",
"10001000111",
"10000010000",
"10000011010",
"10000100000",
"10000001110",
"10000100010",
"10000010011",
"10000011110",
"10000011111",
"10000111111",
"10000010101",
"10000001100",
"10000001100",
"10000011000",
"10000111001",
"10001000000",
"10000010011",
"10000100000",
"10000010001",
"10000111100",
"10001000001",
"10000001010",
"10000011100",
"10000010100",
"10000100111",
"10000010000",
"10000001000",
"10001000010",
"10000001001",
"10000010110",
"10000000101",
"10000101111",
"10000000101",
"10000011110",
"10000101100",
"10000001000",
"10000100000",
"10000011110",
"10001001000",
"10001000111",
"10000010001",
"10000010100",
"10000010001",
"10000011011",
"10000001000",
"10000011011",
"10000101001",
"10000001100",
"10000010010",
"10000000110",
"10000100001",
"10000011011",
"10000111101",
"10000000111",
"10000010101",

"01000111111",
"00110011111",
"01001011010",
"01001001111",
"00111000101",
"01001001010",
"01000101100",
"01001001011",
"01000000100",
"01000111111",
"01000011101",
"01000011111",
"01000111010",
"01001010100",
"01001011111",
"00110110001",
"01001011010",
"01001011110",
"01001010001",
"01000110111",
"01000111111",
"01001011010",
"01001011000",
"01001100011",
"01001100011",
"01001011001",
"01000001111",
"01000111101",
"01001000000",
"01001010001",
"01001011010",
"01000001101",
"01000100101",
"01000101011",
"01001000011",
"00111010001",
"01001100000",
"01000110001",
"01001000010",
"01001000111",
"01000010001",
"01000011001",
"01001010110",
"01001000011",
"01001011011",
"01000101010",
"00111100000",
"01001011000",
"01001010000",
"01001010010",
"01000100011",
"01001011011",
"01001100010",
"01000111111",
"01001100001",
"01001010111",
"01000111100",
"00111100001",
"01001011101",
"01001011110",
"01001001000",
"01001010100",
"01001011000",
"01000011101",
"01000101011",
"01001011000",
"01000001101",
"01001001111",
"01001100000",
"01001001001",
"01001100001",
"01001000010",
"01000110111",
"01000101010",
"01001000000",
"01001000110",
"01001001000",
"01000010010",
"01001011010",
"01001000100",
"01001001010",
"00111011110",
"01001001111",
"00101100000",
"01001011010",
"01001011001",
"01001100001",
"00110101100",
"00111001111",
"00110001001",
"01000101101",
"01001011101",
"01001100010",
"01001001011",
"01001100000",
"01001010001",
"01001001110",
"01000010011",
"01001010110",
"01001000010",

"01000010000",
"00101011011",
"01000001000",
"00111100011",
"00100110111",
"01000110010",
"01000010000",
"01001000001",
"00111010111",
"01000100101",
"01000011001",
"00111011001",
"00111011011",
"01001000111",
"00111010000",
"00101001110",
"01000101101",
"01000101011",
"01000110100",
"01000010101",
"01000001110",
"01000011110",
"01000000101",
"01000100011",
"01001001000",
"01001001010",
"00111010111",
"01000110011",
"01000100001",
"00111000010",
"01000101001",
"01000001001",
"01000010101",
"00111011001",
"01000110010",
"00111001110",
"01000101000",
"01000011000",
"01000000110",
"01000111101",
"00111100011",
"00111011101",
"00111010101",
"01000010101",
"01001001100",
"01000001010",
"00110111100",
"01000010111",
"01000100101",
"01000101111",
"01000100001",
"01000101011",
"01001011010",
"00111000001",
"01001001001",
"01000011010",
"01000110000",
"00110001101",
"01000011000",
"01000111000",
"01000001000",
"00110101001",
"01001000000",
"01000010100",
"00111011010",
"01000111110",
"00111010000",
"00111000000",
"01001011000",
"00110111101",
"01000101011",
"01000000001",
"01000001111",
"01000011110",
"01000110001",
"00111011111",
"01000011111",
"00110111001",
"00111010010",
"00111010110",
"01001000110",
"00111011000",
"00111010100",
"00101001000",
"01000101100",
"01000010010",
"01000000110",
"00100101100",
"00111001100",
"00110000111",
"00111011011",
"01000101011",
"00110100110",
"01000000100",
"01000110011",
"01000101011",
"01000110110",
"00111001111",
"01000010010",
"01001000000",

"00111100010",
"00100010000",
"00111010011",
"00101001001",
"00100100111",
"01000001000",
"00110110011",
"01000000110",
"00110000110",
"01000001011",
"00111001001",
"00110011101",
"00111001100",
"01000000000",
"00111001010",
"00100001110",
"01000001100",
"00110001110",
"01000101000",
"01000001110",
"01000001010",
"00100111111",
"00110110011",
"01000010100",
"01000000001",
"00111010001",
"00110011111",
"01000011100",
"00111010101",
"00110100010",
"01000011110",
"00111001001",
"00110010000",
"00101010100",
"01000010010",
"00110111101",
"00111001000",
"01000010001",
"00110010010",
"01000000000",
"00110101000",
"00111000111",
"00100111111",
"00111001111",
"01000101111",
"01000000000",
"00110000001",
"00111000011",
"01000100011",
"01000010110",
"00110011000",
"00110110101",
"01001011001",
"00110110000",
"01001000100",
"00111100000",
"00111001100",
"00100111101",
"01000000001",
"00111010110",
"00110101011",
"00100111011",
"00101011011",
"00110010100",
"00110111100",
"01000000000",
"00101010001",
"00110101101",
"01000101010",
"00110100110",
"01000100010",
"00101010001",
"00110111011",
"01000011001",
"00110101101",
"00110110111",
"00111001101",
"00101001000",
"00111000010",
"00111001000",
"01000110101",
"00111000100",
"00110111000",
"00100100111",
"01000001000",
"00111011100",
"00111011110",
"00011010101",
"00111001000",
"00100111011",
"00111001011",
"01000011111",
"00110100100",
"00111010101",
"01000101110",
"01000010101",
"00111010000",
"00110111000",
"00110000111",
"01000011111",

"00110011010",
"00100001100",
"00110111100",
"00100010110",
"00100100011",
"00111010101",
"00110000100",
"00110101111",
"00101000001",
"00110111100",
"00110011010",
"00100111001",
"00110101110",
"00111000001",
"00101100010",
"00011010111",
"00111010101",
"00110001000",
"00111001111",
"00111011111",
"00101100000",
"00100111100",
"00100110101",
"00100101110",
"00111000001",
"00110110110",
"00110010011",
"00111010101",
"00111010100",
"00110100001",
"01000000110",
"00110110011",
"00110001101",
"00100000111",
"00111001100",
"00110101101",
"00101010011",
"00110011111",
"00101010001",
"00110100101",
"00110011101",
"00110110010",
"00100011101",
"00101000000",
"01000010010",
"00110010011",
"00101011001",
"00110101011",
"00111010101",
"00111000110",
"00110001100",
"00110101110",
"01001010111",
"00110000100",
"01000110010",
"00110011111",
"00110011110",
"00011100001",
"00111001100",
"00110110110",
"00110001001",
"00100111000",
"00101010110",
"00101010110",
"00110110110",
"00111100001",
"00101000101",
"00100111110",
"01000010101",
"00110010010",
"00110100010",
"00100110111",
"00110101000",
"00110111101",
"00110100111",
"00110110101",
"00100110000",
"00011011001",
"00101001110",
"00110110001",
"01000001111",
"00110011000",
"00101010100",
"00001010011",
"00100101100",
"00101001100",
"00110100010",
"00010100011",
"00101100000",
"00011010111",
"00110100010",
"00111011111",
"00101001101",
"00101001101",
"01000100001",
"00110110100",
"00101001111",
"00110100101",
"00110000100",
"00111001001",

"00011010010",
"00011000011",
"00110100100",
"00010110111",
"00100010001",
"00111001110",
"00101010101",
"00010001011",
"00100101111",
"00110110000",
"00110011001",
"00100110110",
"00110101010",
"00110011000",
"00101100000",
"00010110110",
"00101001110",
"00101011111",
"00110001110",
"00101010100",
"00100100001",
"00100110110",
"00100100010",
"00011000100",
"00110111110",
"00110001101",
"00101010100",
"00111000111",
"00110010100",
"00100010000",
"00111011100",
"00110110000",
"00110000011",
"00010110011",
"00110101110",
"00100100111",
"00100111000",
"00100110110",
"00101001101",
"00101011001",
"00110011011",
"00110010101",
"00010111100",
"00100111111",
"00111010101",
"00100011001",
"00100110110",
"00110000111",
"00110110001",
"00110111010",
"00110000010",
"00110010010",
"01000111110",
"00100110011",
"01000010101",
"00100100100",
"00110000110",
"00011011101",
"00100001001",
"00110010110",
"00101100011",
"00011001011",
"00101000000",
"00101010010",
"00100101011",
"00110110010",
"00100111011",
"00100001111",
"00111000011",
"00110010000",
"00100110000",
"00100110011",
"00110100100",
"00110110000",
"00100101100",
"00110100100",
"00100010000",
"00001000111",
"00100100110",
"00100111000",
"00110000110",
"00100010101",
"00101010010",
"00000111010",
"00100010010",
"00100101101",
"00100100000",
"00010100010",
"00011100011",
"00011000101",
"00110001010",
"00111011100",
"00100111111",
"00100100001",
"00110000101",
"00110000111",
"00101000011",
"00110100000",
"00101011101",
"00101011111",

"00010101110",
"00010110110",
"00101000010",
"00010110000",
"00100000100",
"00101100011",
"00100010110",
"00010001010",
"00100101001",
"00110101010",
"00100001000",
"00100010010",
"00101100000",
"00101010100",
"00100111001",
"00010001110",
"00011100010",
"00011010000",
"00100001001",
"00011010000",
"00010111101",
"00100101110",
"00100011011",
"00010001000",
"00011001101",
"00110000001",
"00101001100",
"00101001101",
"00110000010",
"00100000101",
"00110110101",
"00110100010",
"00100110000",
"00010001000",
"00110100110",
"00100001010",
"00100100101",
"00100000111",
"00100111110",
"00100000011",
"00110001011",
"00101001000",
"00010101010",
"00100110010",
"00100110011",
"00010111110",
"00010100111",
"00110000001",
"00110101101",
"00101001101",
"00101001101",
"00110000001",
"01000101001",
"00011011001",
"01000001101",
"00100100010",
"00110000011",
"00011010110",
"00010101010",
"00100010101",
"00100111010",
"00010101011",
"00011010101",
"00010010010",
"00011001011",
"00101001111",
"00010100100",
"00100001110",
"00110101111",
"00011001010",
"00100101000",
"00100101101",
"00110001111",
"00110100000",
"00100100100",
"00110100001",
"00011100001",
"00000111001",
"00100010101",
"00011011100",
"00101100000",
"00011100001",
"00101001111",
"00000101110",
"00100000000",
"00010111011",
"00000111011",
"00010100001",
"00010011100",
"00010111100",
"00011010011",
"00100010111",
"00011010011",
"00100010110",
"00101001011",
"00101100000",
"00100010011",
"00110001010",
"00100110111",
"00100111010",

"00010000001",
"00010110000",
"00011010111",
"00010100100",
"00011000001",
"00100100100",
"00010011001",
"00010000111",
"00100101000",
"00110001101",
"00001000011",
"00011001001",
"00101000100",
"00100011111",
"00100000101",
"00001100011",
"00011011000",
"00010001100",
"00100000110",
"00011000110",
"00010100110",
"00100100011",
"00100000110",
"00001000101",
"00010100000",
"00011001110",
"00101001000",
"00100111111",
"00101011011",
"00011001001",
"00110101111",
"00101011001",
"00010010111",
"00001000101",
"00101001010",
"00011100011",
"00010100011",
"00010111110",
"00100101111",
"00010101001",
"00100001111",
"00100111111",
"00010011101",
"00100000111",
"00100101001",
"00010100100",
"00010011111",
"00101000101",
"00100100100",
"00010110110",
"00100101010",
"00100001110",
"00111000111",
"00011001100",
"00100011001",
"00011011111",
"00011011100",
"00010110010",
"00010011111",
"00011000001",
"00011010001",
"00010010111",
"00010001000",
"00001011001",
"00010111000",
"00011000110",
"00010010101",
"00100001010",
"00011011101",
"00011000001",
"00010101110",
"00010110001",
"00110000110",
"00110010010",
"00100010100",
"00101100001",
"00011011001",
"00000110110",
"00011100010",
"00011011010",
"00011010000",
"00010101110",
"00100000110",
"00000101101",
"00001000110",
"00010011001",
"00000100011",
"00010100000",
"00001011001",
"00001010010",
"00011001100",
"00011011011",
"00011010000",
"00011001101",
"00101000001",
"00101010111",
"00011011001",
"00100111111",
"00011011100",
"00100100011",

"00001000111",
"00010001010",
"00011000111",
"00010011101",
"00010111100",
"00011100000",
"00010000001",
"00001011111",
"00100000010",
"00101000010",
"00000110100",
"00010001011",
"00000111100",
"00010101100",
"00010111101",
"00001000101",
"00011010100",
"00010000110",
"00010101010",
"00001001110",
"00010011010",
"00100010111",
"00010101010",
"00000100001",
"00000011110",
"00010101111",
"00100001101",
"00010111110",
"00100110010",
"00010110100",
"00100110000",
"00101000001",
"00001000000",
"00000011010",
"00000100101",
"00010111111",
"00010010100",
"00000101001",
"00100100010",
"00001001100",
"00100001000",
"00100111010",
"00010010000",
"00010000111",
"00100001001",
"00001000100",
"00001011000",
"00100100100",
"00011000001",
"00010011100",
"00011001010",
"00010001110",
"00100101001",
"00010110010",
"00011011011",
"00011000001",
"00011011001",
"00010010001",
"00001011010",
"00010100011",
"00000001110",
"00010010011",
"00001010011",
"00001001100",
"00010100001",
"00010010001",
"00010000100",
"00011001001",
"00011010110",
"00001011010",
"00000111010",
"00000011001",
"00100001000",
"00101000100",
"00100000001",
"00100101010",
"00011011000",
"00000101100",
"00010110010",
"00011010100",
"00000111011",
"00010011001",
"00011001010",
"00000100010",
"00001000001",
"00010000001",
"00000100001",
"00010000101",
"00000110001",
"00001001011",
"00010100101",
"00000111010",
"00010110011",
"00001011000",
"00010111101",
"00100100001",
"00011010010",
"00011011000",
"00001011001",
"00100000111",

"00000111000",
"00001011100",
"00010101011",
"00010000000",
"00010100110",
"00011000110",
"00001100001",
"00001000011",
"00010101100",
"00010101101",
"00000011000",
"00000110110",
"00000110110",
"00000000011",
"00010100000",
"00000100011",
"00000110100",
"00001100001",
"00010001010",
"00000110000",
"00001010110",
"00011000100",
"00000011001",
"00000010100",
"00000001001",
"00001011101",
"00011011010",
"00010110111",
"00100000010",
"00001100000",
"00100101011",
"00000110001",
"00000111000",
"00000011001",
"00000011110",
"00010110111",
"00010001010",
"00000100000",
"00100010101",
"00000110101",
"00010111110",
"00100100001",
"00000100010",
"00000101001",
"00010100111",
"00000100100",
"00001010001",
"00001001000",
"00010001000",
"00000110010",
"00011001001",
"00010001011",
"00010110010",
"00000110101",
"00011010111",
"00010100100",
"00010011101",
"00001001100",
"00000111101",
"00001010011",
"00000000011",
"00001000011",
"00001001000",
"00000010010",
"00001001010",
"00001011100",
"00000111001",
"00010001000",
"00001010110",
"00000101101",
"00000011010",
"00000001110",
"00010001101",
"00010111101",
"00011100000",
"00010011111",
"00011000110",
"00000101000",
"00000010001",
"00010111101",
"00000110110",
"00000101101",
"00010001101",
"00000010100",
"00000100100",
"00001100011",
"00000010111",
"00000100000",
"00000010101",
"00000111011",
"00001000110",
"00000001111",
"00010101010",
"00001000011",
"00010100101",
"00010001110",
"00011000110",
"00010100000",
"00001001111",
"00010111111",

"00000101110",
"00000011001",
"00010001100",
"00000000110",
"00000111001",
"00000100000",
"00001010101",
"00000010011",
"00010010011",
"00000000111",
"00000001001",
"00000101110",
"00000010010",
"00000000000",
"00000001101",
"00000011111",
"00000011010",
"00000100100",
"00001100001",
"00000100111",
"00000010010",
"00010010110",
"00000000101",
"00000000111",
"00000000001",
"00000100011",
"00001000000",
"00000010110",
"00001011101",
"00000100101",
"00000010111",
"00000101101",
"00000101101",
"00000001010",
"00000000010",
"00010100100",
"00010000001",
"00000000111",
"00001011011",
"00000101110",
"00010001000",
"00100001111",
"00000011110",
"00000011011",
"00010010100",
"00000100000",
"00000101010",
"00000110000",
"00001001011",
"00000010100",
"00000101011",
"00001100001",
"00010011000",
"00000100101",
"00010001111",
"00001011111",
"00010010001",
"00000110111",
"00000000010",
"00000011110",
"00000000010",
"00000111110",
"00000011110",
"00000000010",
"00000001100",
"00000111101",
"00000011100",
"00001011101",
"00001000101",
"00000011000",
"00000010100",
"00000000111",
"00000101001",
"00000100111",
"00011010011",
"00010000111",
"00000101010",
"00000000001",
"00000001001",
"00010000101",
"00000100110",
"00000100010",
"00001010000",
"00000000011",
"00000011000",
"00000110011",
"00000000111",
"00000010000",
"00000001010",
"00000101110",
"00000001101",
"00000000111",
"00000000101",
"00000100110",
"00000111010",
"00000111010",
"00010000010",
"00010011001",
"00001000110",
"00001001110"


);
end intercon_mem_package;
package body intercon_mem_package is
end intercon_mem_package;
