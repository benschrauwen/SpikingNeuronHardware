library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_signed.all;
use work.settings_package.all;
package weight_mem_package is
constant weight_mem : weight_mem_type := (
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"1011000101001101000011011010100101000110000001100100000000000100001111110101000001011000011100000001",
"0100100001100010101100100100011000000011011110111011000011111100110000010010011110001111000010110010",
"1010101110001110010101010111011100001000111000000111010101111000101000001011010001000100011001111010",
"0011001100101011101010101010100110011000111011001011111001100010000000001011101001110000100101010101",
"0011011100000101000000001110000010100100100010001011010111011101101000101001101111010101011101001000",
"0100000010011001001111000000101011101101100110110011101010100011110110110101011000001101000001110000",

"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"1100100001000000000101000101001101110000100001010010000011010001000000011100100010000000000001100101",
"0011001000111101000010000110110010001100000000101000100110001110100000100010000001011001110000011000",
"0000011010011111100000110001101000101011111010100101100000001011011001011110101100100001010100111100",
"1011110100011100110010000010101100010001111100011110111000101011111110111111001110010100111011111000",
"1010011011001101100100001111101011010110010110100111000000110001111000100110110001011101011100111111",
"0100011100011000001000010010000011010011100110000011110000000010011010010000011010111011011000001001",

"0000100001000001001010000000000000010000001000000001000000100000000000100000001000010000011001000000",
"0000100001000001001010000000000000010000001000000001000000100000000000100000001000010000011001000000",
"0000100001000001001010000000000000010000001000000001000000100000000000100000001000010000011001000000",
"0000100001000001001010000000000000010000001000000001000000100000000000100000001000010000011001000000",
"0000100001000001001010000000000000010000001000000001000000100000000000100000001000010000011001000000",
"0000100001000001001010000000000000010000001000000001000000100000000000100000001000010000011001000000",
"0010101100000011000000000000000000010000011000000011100001110001001000110100001100010010011101001000",
"0001110001111101111111111111001000001101101001100100001110000100010011001011110001001101000000010110",
"1001110111000000001011001111000010110000100101111001111010000100010111001001111011100101111001111001",
"0010001001111101011000100010010110011010001111101001011100010010100010110101000001111001111111010100",
"0111010000011100011011010001110001011110110010010011010010111000001101101101100001010000011101010001",

"0000000000000000000000000000100000000000000000000000000010001000000000000000000000000000000010000000",
"0000000000000000000000000000100000000000000000000000000010001000000000000000000000000000000010000000",
"0000000000000000000000000000100000000000000000000000000010001000000000000000000000000000000010000000",
"0000000000000000000000000000100000000000000000000000000010001000000000000000000000000000000010000000",
"0000000000000000000000000000100000000000000000000000000010001000000000000000000000000000000010000000",
"0000000000000000000000000000100000000000000000000000000010001000000000000000000000000000000010000000",
"0010000000010010000000011000100000001010011000000010100010010000010000000001100000101000110110101010",
"1101110000100001001101100001100101010001000111010000011110001011101111000100011100010010000001010100",
"0010000101001000111011000111100101100111110101111101001000101001111000111110011100000111001010000001",
"0101100011011110110010101000111011000001000100100111101011100100001110101100101111101101001111011111",
"0101011111101001101011010111110000010100001101110011110110011110101001010110000010001001000011100000",

"0000001000100010000000000000010000000000000000011000000000000001000000000000000000000000000000000000",
"0000001000100010000000000000010000000000000000011000000000000001000000000000000000000000000000000000",
"0000001000100010000000000000010000000000000000011000000000000001000000000000000000000000000000000000",
"0000001000100010000000000000010000000000000000011000000000000001000000000000000000000000000000000000",
"0000001000100010000000000000010000000000000000011000000000000001000000000000000000000000000000000000",
"0000001000100010000000000000010000000000000000011000000000000001000000000000000000000000000000000000",
"0010100111000000010011000000010000010000001101011001000110100001000000010000000001001000101100010100",
"1001001000111011101000011111101110100110000010011100011001000101000001101101011000010110010011100010",
"0100001000100110001100101110001011011010110000100110101100000111101100100111000110100000010000100011",
"0010010000110111000110111111110000101001110101011010000000111011001010101000000101100100111011110111",
"1100101101101100110001000100110111101110101100101100001010110110110000011000111111000001110010001001",

"0000000110000010100000000010000000000000000100000000100110000000000011000000001000000000000100001000",
"0000000110000010100000000010000000000000000100000000100110000000000011000000001000000000000100001000",
"0000000110000010100000000010000000000000000100000000100110000000000011000000001000000000000100001000",
"0000000110000010100000000010000000000000000100000000100110000000000011000000001000000000000100001000",
"0000000110000010100000000010000000000000000100000000100110000000000011000000001000000000000100001000",
"0000000110000010100000000010000000000000000100000000100110000000000011000000001000000000000100001000",
"1010000110001010111000010010000000101100000010000000110110010010001111000100101100000000110010000010",
"0001001000110001100100000100001110000010111101101011001100001100100011110011010000011111000100001100",
"0011100011110100000001100010110010010110100100011111000000100101000001001010000100011000000110001111",
"1101111000111011111011111001011100011000010011110110001110100101111011101100100010100001011101011101",
"0100011111100010111001110000011001000001110111111111001101110001010000110010001001110111110000101100",

"0010000001001011001010000000010100000000010000001000000000000000001000001000000100000000100000000010",
"0010000001001011001010000000010100000000010000001000000000000000001000001000000100000000100000000010",
"0010000001001011001010000000010100000000010000001000000000000000001000001000000100000000100000000010",
"0010000001001011001010000000010100000000010000001000000000000000001000001000000100000000100000000010",
"0010000001001011001010000000010100000000010000001000000000000000001000001000000100000000100000000010",
"0010000001001011001010000000010100000000010000001000000000000000001000001000000100000000100000000010",
"0011001001011010001010000100010100010100010000001000000000000000111000100110011110001000100100100000",
"0100000010101101111110110001100010001011101001010011101111001101001011001001100101110011100011011110",
"1100100000100011010011100000010001000000100010001100010011001111001101011000000000001111001000010110",
"0010111101000100111000001101111000100010101010100001101001110011010110011111111011110001110101111110",
"1001111000000011010110011011000011010111100110111010010100110001011000100011111101110110001000101101",

"0000000000000000000000000000000000000010000000000000000000000000000000001110000010000010100000000000",
"0000000000000000000000000000000000000010000000000000000000000000000000001110000010000010100000000000",
"0000000000000000000000000000000000000010000000000000000000000000000000001110000010000010100000000000",
"0000000000000000000000000000000000000010000000000000000000000000000000001110000010000010100000000000",
"0000000000000000000000000000000000000010000000000000000000000000000000001110000010000010100000000000",
"0000000000000000000000000000000000000010000000000000000000000000000000001110000010000010100000000000",
"0001110000010100100010010001000001000010010001110000000001000001010010101010000110000110100100000001",
"0100000111001000010101001100100010110110100100000111001110100110100101010100011010011001111010000100",
"0101001000001011100001000110011100011001001010000110101010000000000101001111101010101111001011001110",
"1110010010111101001101001100000111000000011101000100110000011101111011100000101001000010111011110111",
"1000110101010111000111111000010111111110100011111000000100010101000111000110011110110010011001011010",

"0011000000000001000000000000000100000010100000000000000000000100000000000000000000000000010100000000",
"0011000000000001000000000000000100000010100000000000000000000100000000000000000000000000010100000000",
"0011000000000001000000000000000100000010100000000000000000000100000000000000000000000000010100000000",
"0011000000000001000000000000000100000010100000000000000000000100000000000000000000000000010100000000",
"0011000000000001000000000000000100000010100000000000000000000100000000000000000000000000010100000000",
"0011000000000001000000000000000100000010100000000000000000000100000000000000000000000000010100000000",
"0011000010100111110101001000010100000011010000100101001011110101000000001000001100011110000111010001",
"1000111000011000000010100101001000111000100111011010010000001000111101110011100011100000111000000110",
"1101010111011001001010000110100011000010100100010010100100000011000111101111110011000000010000000100",
"1101111100000000111100010001001111100110111101000100110111111000011010000111110011000011110000110111",
"1110000001110111100100011101111011011110010000111000011111100000001101010001011110011000000100001010",

"1000000000000000000000000001000100010000000000001000000000000000000000000000000000000000000000000100",
"1000000000000000000000000001000100010000000000001000000000000000000000000000000000000000000000000100",
"1000000000000000000000000001000100010000000000001000000000000000000000000000000000000000000000000100",
"1000000000000000000000000001000100010000000000001000000000000000000000000000000000000000000000000100",
"1000000000000000000000000001000100010000000000001000000000000000000000000000000000000000000000000100",
"1000000000000000000000000001000100010000000000001000000000000000000000000000000000000000000000000100",
"0100001000000100000000001001000101010010111000000010110001000011001010000010010010001010000010010101",
"1010000100011011011010100001000110000100000110111101001010111100010001010100000001110100000100101110",
"1111000110111010001110100111110100001101000010011101000001011000110001110000001100100101011000001110",
"1010100011001011100001110011001010011101101010010000000110000101110111101001101010000000100001001011",
"1010110101110101000100010110011011101010011001101000011000000101011111000001010001001101101110011101",

"0000000000000101000000000000000000000000010000000000000000000000000000000000000000010010000100000100",
"0000000000000101000000000000000000000000010000000000000000000000000000000000000000010010000100000100",
"0000000000000101000000000000000000000000010000000000000000000000000000000000000000010010000100000100",
"0000000000000101000000000000000000000000010000000000000000000000000000000000000000010010000100000100",
"0000000000000101000000000000000000000000010000000000000000000000000000000000000000010010000100000100",
"0000000000000101000000000000000000000000010000000000000000000000000000000000000000010010000100000100",
"0010000110010000100000000000000010000100010001001000000010000000010100001101010010010010110100010110",
"0000010001000111001011001111110101000000000100100100010101110100100011000000101101000101001110101100",
"1001101001101101010101101000000000110001001010100010111000111000111100010000111011110100001010000100",
"0110011000001010101110010110001100110011111000010011100100100001001010110101101000001110100110100011",
"0011000001010111111011011001011001111010010000010100001000011011100010011111101100001101010101010110",

"0000010001000000000010001000000000000000000000000000000000000000000000000000000010000000000010000001",
"0000010001000000000010001000000000000000000000000000000000000000000000000000000010000000000010000001",
"0000010001000000000010001000000000000000000000000000000000000000000000000000000010000000000010000001",
"0000010001000000000010001000000000000000000000000000000000000000000000000000000010000000000010000001",
"0000010001000000000010001000000000000000000000000000000000000000000000000000000010000000000010000001",
"0000010001000000000010001000000000000000000000000000000000000000000000000000000010000000000010000001",
"0000110101001001000010001010010111001000010000011000100010001110010000100000001000100011010010000001",
"1001001000110100101111111100101000000000100100000101011100110001101011010110000111011100100001011010",
"1100110011010100011011100000001100000001001101100100000000100000001101111011000110010000100110010110",
"0010001101010011110110001001110000010011111111101110100101100001111101001111101100001110001001100111",
"1011001010011011010000100010001000110100010000111010110101001110010100001100111101001001100010001110",


"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"1101001000001100110010001000000011000100000100000001001000000001100001001011000000101001011100001000",
"0000000010000010001001010110100000011011100000000100010001011010001110110001010001010110100011110010",
"0111001010001101110110111000100100010001110011111011000000110010001101100110101010000111011111111101",
"0000111111000100000011010010110010101110001111111010110100000000110100011110001100110010010110011110",
"0100110010111101100111000110011111101011111101011100011111000111010100011110101011000011001101000100",
"0000100001010001001011110111111011111011101101100011001110000110000101001010001011010011011110010001",

"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"0111110001011000001001000100010001100100101101010000101010110010000000010100010001100000011110111001",
"0100000100000101000000010011101100010001110010100101011101001001101000100011101000011010001000010011",
"0000010111000110101110010111011100001111010111111001010011010010101001011011110100001011100110000110",
"1010111111000011010110101111000110011001010001111101110001001100011111010010110111010111110010000100",
"1001010101100110111111101010010111110010000000001001100000100011111110001000101000100100100110100100",
"0000110010010001011111001111101001110110011111101010001110000101010110110011001100110010110101000011",

"1000000000000000000100000010000000000010010000000000000000000000000000010000100000000001010100000000",
"1000000000000000000100000010000000000010010000000000000000000000000000010000100000000001010100000000",
"1000000000000000000100000010000000000010010000000000000000000000000000010000100000000001010100000000",
"1000000000000000000100000010000000000010010000000000000000000000000000010000100000000001010100000000",
"1000000000000000000100000010000000000010010000000000000000000000000000010000100000000001010100000000",
"1000000000000000000100000010000000000010010000000000000000000000000000010000100000000001010100000000",
"1000011010010000000100100010000100100110001000010001000010000000010000010101100000000001001101110000",
"0101100000101101110101001001110010011000110111001010101001100011000111101000010100110111110000001111",
"0100100001001000010100001101101011100010010110100000100001111101001010101010110100000001110100000000",
"0100011101111111001010000100001011000010100100000111010001100101011100010011100010101101011111101110",
"0011101010110011011110010110010010000111111010100111010100100001100010100100001101000101000111100110",

"0000000000000001100000000100000000001000000000000010000010000000000000000000000000001000000000000001",
"0000000000000001100000000100000000001000000000000010000010000000000000000000000000001000000000000001",
"0000000000000001100000000100000000001000000000000010000010000000000000000000000000001000000000000001",
"0000000000000001100000000100000000001000000000000010000010000000000000000000000000001000000000000001",
"0000000000000001100000000100000000001000000000000010000010000000000000000000000000001000000000000001",
"0000000000000001100000000100000000001000000000000010000010000000000000000000000000001000000000000001",
"0010001001000001110001000100000000101010001011101010101110000000000110010000110001010000101100100001",
"0100010000110101100100000001100110010001100000010010000010100010010001100000000010101001010010000110",
"1001010100110100100110010111110111010101010100000000010100000100101001100111001110001011100011001010",
"0100110010011111111100101011011100011001001101100100100011111101110010111011111111111111001111111001",
"0011001100101101111100000110100010100000010001000001110011001011110011010011101010100000011010110101",

"0000000110000000000000000000000010110000000000000000000000001000000000000000001100000001000001001001",
"0000000110000000000000000000000010110000000000000000000000001000000000000000001100000001000001001001",
"0000000110000000000000000000000010110000000000000000000000001000000000000000001100000001000001001001",
"0000000110000000000000000000000010110000000000000000000000001000000000000000001100000001000001001001",
"0000000110000000000000000000000010110000000000000000000000001000000000000000001100000001000001001001",
"0000000110000000000000000000000010110000000000000000000000001000000000000000001100000001000001001001",
"0000001110000000000000000000000000110001010000001100000000000001001010010000001000100101001001001011",
"1000110100110010110011100110000011001000000011100011010111111110010001000111011100010010100111001001",
"1111010001001100011100000111011111110110101110000000101111011100100000101101011101000011010111100000",
"1000011010011101001110011010100011010111000001111001111101100011110100001111101011001010111100111101",
"1010111100111100001010110110010001111111001000001110001001111100010110000110100011010010111110101110",

"0000000000001000001000000000100010000100000001000000000000000011000000000100010000000000000000000000",
"0000000000001000001000000000100010000100000001000000000000000011000000000100010000000000000000000000",
"0000000000001000001000000000100010000100000001000000000000000011000000000100010000000000000000000000",
"0000000000001000001000000000100010000100000001000000000000000011000000000100010000000000000000000000",
"0000000000001000001000000000100010000100000001000000000000000011000000000100010000000000000000000000",
"0000000000001000001000000000100010000100000001000000000000000011000000000100010000000000000000000000",
"0000000000001010001000110010100010001110000001000100000000010011100100010100011000000010010101000111",
"0001001101101000100111000101011111100001110100000011100001101101010011101011000010110101000010011000",
"1100011000110001011110000100111110100000110010110100010010100110011110001001010110111001101001001001",
"0011110010000110000100001011110100110110001010001001110110010010100001010001101001001110100010110000",
"1011110111001111010011010100001111011110001111100001101001010101011000000010010111011110110010010000",

"0000000001010000000000000000000000001001001000010000000001000001001000000000001000110000000000100000",
"0000000001010000000000000000000000001001001000010000000001000001001000000000001000110000000000100000",
"0000000001010000000000000000000000001001001000010000000001000001001000000000001000110000000000100000",
"0000000001010000000000000000000000001001001000010000000001000001001000000000001000110000000000100000",
"0000000001010000000000000000000000001001001000010000000001000001001000000000001000110000000000100000",
"0000000001010000000000000000000000001001001000010000000001000001001000000000001000110000000000100000",
"0000010011010010000010000010000001001001011010011011010101010101011001000000000000101010100000010000",
"1111001000001101110100100101111100110100100001100000100011001001001000011011011001110101011110101101",
"0111001101111000111001001000110000110001100010000000100011100000100010111011111010010001000011100110",
"1011111100111100010011110100010010111110010000100101011100111000001100000101111001010000101010011111",
"0110010001110001100010110010100101110000100101011111110001101011011001001000001101100110010001011101",

"0000000101010000000000000000000001000000000001000000000000000000010000000000010000000000001000000000",
"0000000101010000000000000000000001000000000001000000000000000000010000000000010000000000001000000000",
"0000000101010000000000000000000001000000000001000000000000000000010000000000010000000000001000000000",
"0000000101010000000000000000000001000000000001000000000000000000010000000000010000000000001000000000",
"0000000101010000000000000000000001000000000001000000000000000000010000000000010000000000001000000000",
"0000000101010000000000000000000001000000000001000000000000000000010000000000010000000000001000000000",
"0010100111110000100100100000000101001000100011001000010001100001010000000000010000110100001010010001",
"1001011000001010011000000111101000000111010101010110001000010100011001101011100111001011100000101110",
"1100011001000100000011000111110010010111000101100001001110000110110001110011011000001110010001100100",
"0011010010100011101100101101000111110100011010100111010110001000100110010011100111010010100111011000",
"1010010001011111000101011101110110100011001111001101101000000100111100101110000101000011100011111111",

"0000000000000000000010000000000000000000100000000010000000000000100000000000000000000001000000110000",
"0000000000000000000010000000000000000000100000000010000000000000100000000000000000000001000000110000",
"0000000000000000000010000000000000000000100000000010000000000000100000000000000000000001000000110000",
"0000000000000000000010000000000000000000100000000010000000000000100000000000000000000001000000110000",
"0000000000000000000010000000000000000000100000000010000000000000100000000000000000000001000000110000",
"0000000000000000000010000000000000000000100000000010000000000000100000000000000000000001000000110000",
"1000000010000000000011100000001000010010100000001110101001000100110001000101000000000010010001110000",
"0100111100010000111110011111010100100101011111110010000100010001101000111010000111000101001000110011",
"0111101100101110101110010010000011101001110101011001110010000010110100101010110001011001100100000111",
"1011010010001111100001100100111000110000011100110110010100110111101010111101111010110111000110011101",
"1011010001000111111111011011001001101011111101110101000101101110001100111110010101000001111100011010",

"0000000000000010000000000010001000100000000000000000010000000100000000000100000000000000000000000000",
"0000000000000010000000000010001000100000000000000000010000000100000000000100000000000000000000000000",
"0000000000000010000000000010001000100000000000000000010000000100000000000100000000000000000000000000",
"0000000000000010000000000010001000100000000000000000010000000100000000000100000000000000000000000000",
"0000000000000010000000000010001000100000000000000000010000000100000000000100000000000000000000000000",
"0000000000000010000000000010001000100000000000000000010000000100000000000100000000000000000000000000",
"0100001101100110010010010110101010100000000001000000100100000110010000110111010011001000000011000000",
"1000110010001011001101101011011000111100111100111101010001110101001100001000101100110011010100101101",
"1001110000010000110000001010001101101011011010001111011001001100100111101100000100000011110000111110",
"0110100110001101101111011010101111101000000001111110110011100001010100000011010110000100101011001101",
"0110011011001001100100101100110011011100100101101111010011101010100110010010001110011100010110101000",

"0000000000001000000000000000010000000000100000000000000000000000000001000010000000100000011000000000",
"0000000000001000000000000000010000000000100000000000000000000000000001000010000000100000011000000000",
"0000000000001000000000000000010000000000100000000000000000000000000001000010000000100000011000000000",
"0000000000001000000000000000010000000000100000000000000000000000000001000010000000100000011000000000",
"0000000000001000000000000000010000000000100000000000000000000000000001000010000000100000011000000000",
"0000000000001000000000000000010000000000100000000000000000000000000001000010000000100000011000000000",
"1100000000001010100010000100010010011110100000100000000011000000100001100010100000000000011001000000",
"0010001011001101001000101001101100000001010001010110011000001111001011011101000110100010000010010010",
"1001011100011001011100100110100101100011100111010111011000101100011101011111011011111101010010101111",
"0001110011111111100111011011110010100100011111111100001110011001010010001000111111000011100100000111",
"0110100101000000101101000000010011101100001100000011101110001101111110111101110101101100110000101011",

"0000000000000000000000000000000000000011000000000001000000000010000010000000000000010000000000010000",
"0000000000000000000000000000000000000011000000000001000000000010000010000000000000010000000000010000",
"0000000000000000000000000000000000000011000000000001000000000010000010000000000000010000000000010000",
"0000000000000000000000000000000000000011000000000001000000000010000010000000000000010000000000010000",
"0000000000000000000000000000000000000011000000000001000000000010000010000000000000010000000000010000",
"0000000000000000000000000000000000000011000000000001000000000010000010000000000000010000000000010000",
"0100010000000000101001000010000000001101001000000001010000000010010010000000010000010000100010010000",
"1010100010011001000100111100100101000011010101111001001111101001101101011001100100100110001100100111",
"1011000111001111000010010101101101110011111001011000101111101101001001010000000111111111110000000011",
"1011101001111100011111110000010010001100010011000110011101010111001101100011101100111001010101101011",
"1010111111101100111000100101110001011010010010001111101000011111011001110111101110011010000011110010",


"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"0110110111000100010001100010100000010000000101001010101000101000011011010110010111110100110110101001",
"0001000000110001101101011110001111101011011011110000010100100111000000110000001000000001000000000010",
"0110111010110000111010111101111001110101100110011001100111001110010110001000100101111001110110010010",
"0100101001000000000100010100100101111010010110101111011000011111110100101101110011111010100111110100",
"1011111101101110101100100100111000000110001010110001100010000000011011101110111010101000001101100100",
"0101000000110101111011101000110101000111000110111010100010000110110100011011010001101110010100011110",

"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"1000000010101100101010000101100111101100111101010001011010100000010100000010100100001000101001010000",
"0000111000100110010001110000000000000000100010011100100101010110001010111000110011010111000000001100",
"1010111110010011111000011111111010010100001100100110110000111100110000100110010100010011101101110010",
"1011111101011000001001100000011101110100001011000000010000000001101011110011001011110011000100100010",
"1110110111011001101111000000110100010011000000001110100001101000110001101101001111001111110110101011",
"0101111001010001100100010110110001001110100110010111010001011000011001101011011100110110000101010010",

"0000000100100000000000010100000000101000000000000000000000000011000000001000000000000000001000010010",
"0000000100100000000000010100000000101000000000000000000000000011000000001000000000000000001000010010",
"0000000100100000000000010100000000101000000000000000000000000011000000001000000000000000001000010010",
"0000000100100000000000010100000000101000000000000000000000000011000000001000000000000000001000010010",
"0000000100100000000000010100000000101000000000000000000000000011000000001000000000000000001000010010",
"0000000100100000000000010100000000101000000000000000000000000011000000001000000000000000001000010010",
"1011000110000100100010011100000000101000100100000000000100010110000101001110100000000110001000010110",
"0100110000110000011100100100111001101101001000001111011000000011011010110000000010100000111111010011",
"0010010000100011100101010001010111010100011000110101110001010001110010100100010001101011101110101001",
"1001011111111011010101111011011001000010010110111101001011101110000000000010101000001000001111111100",
"0001110010010110011000100101011111001100001101111000101100001011110000001001010100110000011000110111",

"0000000000000000010000000000000110000000001000001000000000000000000010000000100000010010000000000011",
"0000000000000000010000000000000110000000001000001000000000000000000010000000100000010010000000000011",
"0000000000000000010000000000000110000000001000001000000000000000000010000000100000010010000000000011",
"0000000000000000010000000000000110000000001000001000000000000000000010000000100000010010000000000011",
"0000000000000000010000000000000110000000001000001000000000000000000010000000100000010010000000000011",
"0000000000000000010000000000000110000000001000001000000000000000000010000000100000010010000000000011",
"1100101011000100110100011010001110010000001000001000000001010011100111000010101001011010000000001011",
"0011000000010000010011000000010001100100110010101101001010101000010000001101110010100010100011110110",
"0011010000010010000000100100010111100011111001010101101100001100011110111000110100010100100101100001",
"0101101110101111111110011111111110001000101100110010110101010000011001101101100110111001111011111111",
"1100111101101101000010011110011001111111111100101011010111100001001000100110011010000111000010000101",

"0000000000000000000000000000000000000010000000000000000011000000000000100010010000000010000000000000",
"0000000000000000000000000000000000000010000000000000000011000000000000100010010000000010000000000000",
"0000000000000000000000000000000000000010000000000000000011000000000000100010010000000010000000000000",
"0000000000000000000000000000000000000010000000000000000011000000000000100010010000000010000000000000",
"0000000000000000000000000000000000000010000000000000000011000000000000100010010000000010000000000000",
"0000000000000000000000000000000000000010000000000000000011000000000000100010010000000010000000000000",
"1100011000100010000000000010000011101110000000000010010011100010000001100111010110010110000000000001",
"0001000011000100101100110001111000010001110100100100000011010000101010000010010001100010010111111000",
"0000010111011000001001001101100100010001010001011011101100000001111100110000111001101011111011101010",
"1000101001111101100110000010101101100110010110111100001111001100110101111111101101011101101011001101",
"0111100011001010011000011110111111001001101001000100101000101011010101110100000100011100010100000000",

"0000001000100000000000000000001010010010000000000010000000000100000000000000000000000000000000000100",
"0000001000100000000000000000001010010010000000000010000000000100000000000000000000000000000000000100",
"0000001000100000000000000000001010010010000000000010000000000100000000000000000000000000000000000100",
"0000001000100000000000000000001010010010000000000010000000000100000000000000000000000000000000000100",
"0000001000100000000000000000001010010010000000000010000000000100000000000000000000000000000000000100",
"0000001000100000000000000000001010010010000000000010000000000100000000000000000000000000000000000100",
"1110001000101000000000001110100010110110001000001001000100000101100000000001000001001000000110001011",
"0001111011010100001101100001011111011001110111100110100010001000001001001110011010010111101001110100",
"0001101111110111110110110000011101001010010111110010100011110100000111100000111010110000110101001100",
"1010101110011111010110101111110000000001110000101001111100000000010111011111100101101101001001100111",
"1001011000001100000001001000111110011011110111111010101111101111000110011010101010111110011011100101",

"0000000000001100000010000000000100010000101100100000000001000100000000010100010000000000000000100000",
"0000000000001100000010000000000100010000101100100000000001000100000000010100010000000000000000100000",
"0000000000001100000010000000000100010000101100100000000001000100000000010100010000000000000000100000",
"0000000000001100000010000000000100010000101100100000000001000100000000010100010000000000000000100000",
"0000000000001100000010000000000100010000101100100000000001000100000000010100010000000000000000100000",
"0000000000001100000010000000000100010000101100100000000001000100000000010100010000000000000000100000",
"0010000000001110001010000000001100000010111000001001100001010100000000011100110000100000000000000001",
"1101111111000001100100001011110010010101001111110010001111001000011101000111001110011111000011100100",
"1101101000010001100110110100000110111100000111100000010111100011011111000110011010000011111110111010",
"1010110100101011010001101100011111111111010110000111101011000011100000101011111101000010010100100101",
"1101100010011011110100101000101110100001010000111101101110100111010100010100110000110011100001010100",

"0000000000000000000000000000100000000000000001100000000000000000001000000000000000000000000000000000",
"0000000000000000000000000000100000000000000001100000000000000000001000000000000000000000000000000000",
"0000000000000000000000000000100000000000000001100000000000000000001000000000000000000000000000000000",
"0000000000000000000000000000100000000000000001100000000000000000001000000000000000000000000000000000",
"0000000000000000000000000000100000000000000001100000000000000000001000000000000000000000000000000000",
"0000000000000000000000000000100000000000000001100000000000000000001000000000000000000000000000000000",
"0000000101100001000000100000000000010000001001100101100000000000000000000011010000010100100001100010",
"0111011010001000011110010101100101101101010101100000011000111011001100010000101001101011000000011001",
"0011110000001110101001010111111010001100100000001000000111101011111101001100001101101111001100011101",
"1100111001111101100110000111100110000111100010111001110100011001101010100100010001010010110110100101",
"1110010100000111010101011000110101101100101011010010100001111110010001111111110111100011100001100110",

"0000000000000000000000000000000000000000000000000010000000000000000000000000010000000001000000000000",
"0000000000000000000000000000000000000000000000000010000000000000000000000000010000000001000000000000",
"0000000000000000000000000000000000000000000000000010000000000000000000000000010000000001000000000000",
"0000000000000000000000000000000000000000000000000010000000000000000000000000010000000001000000000000",
"0000000000000000000000000000000000000000000000000010000000000000000000000000010000000001000000000000",
"0000000000000000000000000000000000000000000000000010000000000000000000000000010000000001000000000000",
"1000000010010100000000101010101000001000001000100100011000000000000000111100110011000001010000000000",
"0110110101100011001100010100010011010101110011011010100001110101011110000000011100011011101110101010",
"0001111101001011010101110000010000110101000100000010010011110101001111000001001000000001100001110110",
"0111000101110001011010011101100110011011110001000100100110011010100111001110101010111100111010101111",
"1100110100001001110100001100111011111011000011001101101100010011110001001001001110001001001111000111",

"0100010000100100000000000010000110011000000100010000000001000000011010000000000000110000001000000000",
"0100010000100100000000000010000110011000000100010000000001000000011010000000000000110000001000000000",
"0100010000100100000000000010000110011000000100010000000001000000011010000000000000110000001000000000",
"0100010000100100000000000010000110011000000100010000000001000000011010000000000000110000001000000000",
"0100010000100100000000000010000110011000000100010000000001000000011010000000000000110000001000000000",
"0100010000100100000000000010000110011000000100010000000001000000011010000000000000110000001000000000",
"0110010000100100001000000010100110010010110100010000000001100000011010000011010000110101000000001100",
"1000101011001101110001001110011010001001000101110110001000011111000011111000101001111010001101110010",
"1111110111101000000110011010111010101000001001111100110111101010110111011100101011000000111100110001",
"1101011110011011001100100100000101011110011011000101001111011011110110100111011101001000011110101110",
"1001110010010110011000010001010001110011001100011000110101001111001100011000001110100100101100001000",

"1011000000100000010000001000000010010000100000001010000000100000000101100011110011010001000000110000",
"1011000000100000010000001000000010010000100000001010000000100000000101100011110011010001000000110000",
"1011000000100000010000001000000010010000100000001010000000100000000101100011110011010001000000110000",
"1011000000100000010000001000000010010000100000001010000000100000000101100011110011010001000000110000",
"1011000000100000010000001000000010010000100000001010000000100000000101100011110011010001000000110000",
"1011000000100000010000001000000010010000100000001010000000100000000101100011110011010001000000110000",
"1111000001100000011000100101000110000000100000110010000010000000010010100010110011110001000000110110",
"0000001000000001100100001000111001011110110011001010000001110101001101100001001000011101110011001000",
"0001110110110011010111011011001011010111111100001111110001101010001101111011000010000010011000010101",
"1000000101111110111110011100110000100101000011101110101110011111110011111000000101111101100011100001",
"1011110111100100101110101010111010101001101101110000111011100011110111100110011010001011001111010010",

"0001010000001100010000101000001000000000000000000000000000000000000000000100000000000001010000000000",
"0001010000001100010000101000001000000000000000000000000000000000000000000100000000000001010000000000",
"0001010000001100010000101000001000000000000000000000000000000000000000000100000000000001010000000000",
"0001010000001100010000101000001000000000000000000000000000000000000000000100000000000001010000000000",
"0001010000001100010000101000001000000000000000000000000000000000000000000100000000000001010000000000",
"0001010000001100010000101000001000000000000000000000000000000000000000000100000000000001010000000000",
"0101110101001100010010111000011100010000000000000000100000010101011000001000101011100011110000000100",
"0011010000011110100000101011001000101001001110101100001110100000000101000111010000010101011001111001",
"1010001010001001001101000110100011000100110011110101000101000101001100111101010100000001111011000000",
"0000001010111011000101010001000000011000001111101000010010011010100111000100101010011101000111110111",
"0100100011100111111000100011100110100011000100001010111101010000100011000010000000101011011110001101",


"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"0111001011101000111100010110110100110111000011100001111000000111101101010101111111100000000001000100",
"1010000100000101000011001001000010001000110010000110000110111000000010101000000000011011011101000011",
"0000011000110111101011000110111001101010110001001101101110101110110001000110011100000110100110011100",
"1001111010101101111111111100011010100010011100110100101010100000101000100000001101111000010000111001",
"1101001100011011100100001010010101111001000100000111011001000110111000010100010111010011000000001111",
"1111011001001011100100100111110101110100110010001001100010110111011111110000001110001010011011001010",

"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"0111010011001110000100101000000111010110001000000010111000111010011000010000010110010011101001110111",
"0000101100100000100010001000001000000101010100100101001000010001001100000111001101000001010011000000",
"1110101100100010110111110111111110001011010111011101010110000101000101111101010001100010110100111001",
"0110001011111001001100010110011111100011100101110100010111101011010110111000010011100010011100100001",
"0001101100010011010011001011000000100001011110000000010011101001101011000111110000111100011001011000",
"0010010101010011001110110010011011010000001000100110001111110001010100010111011011000000100110000001",

"0000010000000101000000000000001001000000000010001001100000010000000000000010000000000001000000000000",
"0000010000000101000000000000001001000000000010001001100000010000000000000010000000000001000000000000",
"0000010000000101000000000000001001000000000010001001100000010000000000000010000000000001000000000000",
"0000010000000101000000000000001001000000000010001001100000010000000000000010000000000001000000000000",
"0000010000000101000000000000001001000000000010001001100000010000000000000010000000000001000000000000",
"0000010000000101000000000000001001000000000010001001100000010000000000000010000000000001000000000000",
"0100010010000000001000001000011001000010000011001001111100010000000000000111000010000001000011010000",
"0010111100110101100001100001000000000101001000001001000011111010001111010000110001111100001100000110",
"1001010001010101010000110010110111111101110100111110000010110111100010110000010000001000011000001111",
"1010100100011011011110000101000011000100111001100101111011000101010111001101011101100100100010111100",
"1001111001011100010101111101100110011100011110011010101110111011101111000101111001110111011001111101",

"0000100000000000000000000000000000001000000000000000000001000000000000000000000000010000000100100000",
"0000100000000000000000000000000000001000000000000000000001000000000000000000000000010000000100100000",
"0000100000000000000000000000000000001000000000000000000001000000000000000000000000010000000100100000",
"0000100000000000000000000000000000001000000000000000000001000000000000000000000000010000000100100000",
"0000100000000000000000000000000000001000000000000000000001000000000000000000000000010000000100100000",
"0000100000000000000000000000000000001000000000000000000001000000000000000000000000010000000100100000",
"0000100010001000001000000101000100001010000100000000001001010000000000000000000110010011000110100100",
"1010001000110010000001011010110000111001100010101101110111100010111101100111111000011100100000000000",
"1111011010000101100101011010101100100100010011100010101011011101001111010010101000100101111101110010",
"0110011100001010110000111010111011101000110000011001100000001110010100111000010101011010000000111101",
"1001100101101010000011000110100010001111011101011111110110100101010011101001101000100010010111100010",

"0000100100000000000000100000000000000100000000000001000000000000010000000000001000000000000001000000",
"0000100100000000000000100000000000000100000000000001000000000000010000000000001000000000000001000000",
"0000100100000000000000100000000000000100000000000001000000000000010000000000001000000000000001000000",
"0000100100000000000000100000000000000100000000000001000000000000010000000000001000000000000001000000",
"0000100100000000000000100000000000000100000000000001000000000000010000000000001000000000000001000000",
"0000100100000000000000100000000000000100000000000001000000000000010000000000001000000000000001000000",
"0011100110000110001000100010000010000100101000100001011001000010111000000100000100000001001101000000",
"1100000001111001100011011001100100101111010101000100100010110100010111011011111010001000010000101011",
"0000011101001000110101101101111001111000010111010100010010111100001000110001011100011110111010000010",
"1000111100011110001011100100000101011100011101111011101100101111100000010110100001111010110001100110",
"1101110000010111000100001100010111101111001010010011000001100000110111101101111000101111010101010111",

"0000000000000000000000000001000100010000100110000000000000000000000000000000000000000000000100100100",
"0000000000000000000000000001000100010000100110000000000000000000000000000000000000000000000100100100",
"0000000000000000000000000001000100010000100110000000000000000000000000000000000000000000000100100100",
"0000000000000000000000000001000100010000100110000000000000000000000000000000000000000000000100100100",
"0000000000000000000000000001000100010000100110000000000000000000000000000000000000000000000100100100",
"0000000000000000000000000001000100010000100110000000000000000000000000000000000000000000000100100100",
"1011000000000000001100000001000110010100101111100010010001100000000000000001100110101001111100100111",
"0000001111111111000011001100000001001011010010010001101010010111100000101110011000010110000110010100",
"0100101011110100110001001101001100100011000100000000100100000111111111011110001001000110000000011100",
"1010110011010011111010110111111111001001110110001111111110100001001000010010010011010010010001111001",
"0011001001000010000110000001111101011101111111010111010100101011000111010100001100010111010110101001",

"0000000000000000000100000000000000000010001000000001000000000101000110000000000001000001000010000100",
"0000000000000000000100000000000000000010001000000001000000000101000110000000000001000001000010000100",
"0000000000000000000100000000000000000010001000000001000000000101000110000000000001000001000010000100",
"0000000000000000000100000000000000000010001000000001000000000101000110000000000001000001000010000100",
"0000000000000000000100000000000000000010001000000001000000000101000110000000000001000001000010000100",
"0000000000000000000100000000000000000010001000000001000000000101000110000000000001000001000010000100",
"0110000000101000001111110000011000000010101000000001000110000101100110100001000011000001000111000100",
"1000010110010011000000001101000101010010010111111010001000101000011100000100011000011100011010101100",
"1000110001000001100000000110000011011011001111000111101011111011010011000100100100010011111010110010",
"0011101110001001111000010101100111110100101110010100101101000001001100011000111111100000011101001111",
"1110010111010110100100110001000000110100110111111011110101110010100011100111000100011111001111101111",

"1000000000000000001000000000000100000100000000100000000011000100000001010000010000001000000000010000",
"1000000000000000001000000000000100000100000000100000000011000100000001010000010000001000000000010000",
"1000000000000000001000000000000100000100000000100000000011000100000001010000010000001000000000010000",
"1000000000000000001000000000000100000100000000100000000011000100000001010000010000001000000000010000",
"1000000000000000001000000000000100000100000000100000000011000100000001010000010000001000000000010000",
"1000000000000000001000000000000100000100000000100000000011000100000001010000010000001000000000010000",
"1000001001000000001100111010100100001100001000101010000101000100100101010110111010001011000001010000",
"1110000010110111100000000000011000100100100101010100111010010010011011001001010001010100101000100011",
"0111110010100100011001000001001110000110000000000000011010000001011000111001001010111000100110111110",
"1111100110101010010110010000110010011011010011000101011110101110111001011110110101110101110011001111",
"0000000110101010011010000110110011110010101011101010101000110100001010001111110001101100010111000111",

"0000010000000100000000000000000100010000000000000000000000000000000001000001100010010001000000000000",
"0000010000000100000000000000000100010000000000000000000000000000000001000001100010010001000000000000",
"0000010000000100000000000000000100010000000000000000000000000000000001000001100010010001000000000000",
"0000010000000100000000000000000100010000000000000000000000000000000001000001100010010001000000000000",
"0000010000000100000000000000000100010000000000000000000000000000000001000001100010010001000000000000",
"0000010000000100000000000000000100010000000000000000000000000000000001000001100010010001000000000000",
"1100000010010101000001011000000111010000000010000001001001000001000001100001100111000001000101100001",
"0000011101001000101000000100010000101001010001100010010010100010111000000110000000110110111010010000",
"1011111100100001100010100100111100110111101101101110010010011110010101110110001110110001111010001100",
"0000011110010100110011000111110000011000010010011001100101111111000100011111011001001100100010001011",
"0110011100011110101100010001000100100001111111001100111101111001111010001000011011110000010110110001",

"1000001000000000010000000001100000000010000000100001010000000000000000100000001000000000000000010000",
"1000001000000000010000000001100000000010000000100001010000000000000000100000001000000000000000010000",
"1000001000000000010000000001100000000010000000100001010000000000000000100000001000000000000000010000",
"1000001000000000010000000001100000000010000000100001010000000000000000100000001000000000000000010000",
"1000001000000000010000000001100000000010000000100001010000000000000000100000001000000000000000010000",
"1000001000000000010000000001100000000010000000100001010000000000000000100000001000000000000000010000",
"0000101010010100010001000001101100000010001010100001010010100111000100000000011010000100000001100000",
"1110010101001000111100111111100001110101100100001001110100010000011001110111101101110000001010010010",
"1010110101101000011110111100000010001011110100011001101011000000101011110100100000011000100000011101",
"1011001000000001100100001000111010101010000101010110111101111101111010001000100111101011100100100000",
"0101000111111111111100110011100001010111011101001001111001110010100101001001101000110001011101100011",

"0000000000000000000000000000000000000000000000000001000000111000000100100000010100000100000000000000",
"0000000000000000000000000000000000000000000000000001000000111000000100100000010100000100000000000000",
"0000000000000000000000000000000000000000000000000001000000111000000100100000010100000100000000000000",
"0000000000000000000000000000000000000000000000000001000000111000000100100000010100000100000000000000",
"0000000000000000000000000000000000000000000000000001000000111000000100100000010100000100000000000000",
"0000000000000000000000000000000000000000000000000001000000111000000100100000010100000100000000000000",
"0000000110000101000000100000101000010100000010000010001001111011100000110000000110100100000100000000",
"1001001001110010110100011111000110100010001101100101000110001100010101101111110001000111010011100110",
"0011100001100010110011011011000101001001111100110101100010101010001111100001111101011111111000100000",
"1101100111111000001110010101011111011110101010101011111111011100111001001111000100011001111011001110",
"1001010010101111100011101110001111100010100100010000000001110001110111010101011011110011100111110101",

"1100000000000100100000000000000000000100000000001000000000000100100000100000000000000001010000000000",
"1100000000000100100000000000000000000100000000001000000000000100100000100000000000000001010000000000",
"1100000000000100100000000000000000000100000000001000000000000100100000100000000000000001010000000000",
"1100000000000100100000000000000000000100000000001000000000000100100000100000000000000001010000000000",
"1100000000000100100000000000000000000100000000001000000000000100100000100000000000000001010000000000",
"1100000000000100100000000000000000000100000000001000000000000100100000100000000000000001010000000000",
"1100000001001110100000000101000011100110000010011100010001000100100101100010001000010001001000001001",
"0101011010100101001100000010111000011100011101000000101010101111010010110101010010100101010101100000",
"0100100100110101111101111110100000011101001000100011100110111001101001001000110111100010110110111010",
"0011110010100000001110001001011010110101100111000101100101011100000010111110110011111001010110100110",
"0000000100110100010011001001000101101010010010100100101110101111000000010100011111011011001001100010",


"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"0110101000000100000110101110100001000100010011001101100001000010000000101010000100000001000010101101",
"0001010011010011110101011000011010100011001000010010000100111001111000000100011010000100111000110000",
"1111010010110100100011010110111010111000010011001100111000001101111010101010001010000011100011011001",
"0000011101011110100011110001000010000100100001101000010111001111011111100000111101011010011111011110",
"1001110111110001001010110100001111011110001100111010010111110110100110001111101101111010000001101010",
"1101111110011000110100100110110100011000001010110000110000110111111000110001101001011111110010010000",

"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"0111101101001000111000101100111110000010001010000101000011011100011010110000111101010010101110000000",
"0111000010100111000001001011000001111001100001110010010000100000010100001100000001011100111100100100",
"1000010010111101110100110011110010010011000000101100100001110011100110101001010100100101000001100111",
"0000100110100010001001100111010111110100111110101111000010001001101101111001000010101001010001001111",
"1000000101110100010110100111001111001010011011110101101101010100100100000011101100001001110001010010",
"0100001011000110000110110110000000101010111111111010011011111001110100101000100000001001011110100000",

"0000000000000001000000000000000000000000001101001000010000000000000011000000001000000000000110000000",
"0000000000000001000000000000000000000000001101001000010000000000000011000000001000000000000110000000",
"0000000000000001000000000000000000000000001101001000010000000000000011000000001000000000000110000000",
"0000000000000001000000000000000000000000001101001000010000000000000011000000001000000000000110000000",
"0000000000000001000000000000000000000000001101001000010000000000000011000000001000000000000110000000",
"0000000000000001000000000000000000000000001101001000010000000000000011000000001000000000000110000000",
"0000001000000011010000000010011001010110011100011010000001000001000011010001110000001100000000100000",
"1001010111001100100101010000000110101001101001101001110100001100001111001010001000110010010110001100",
"0101000010001100001011101101100010101000001101100100011110110011110101101110001111011010111110010111",
"1011100001000000111011001111010110011000110010001101100110111000111001011110011101000001000111001101",
"0000001001110001011000010101000000111000110011011010111101001100010100100100100100110111010100011000",

"0000100000001000000000000000000000010100000000000000110000000001000000000110000000000010001000000100",
"0000100000001000000000000000000000010100000000000000110000000001000000000110000000000010001000000100",
"0000100000001000000000000000000000010100000000000000110000000001000000000110000000000010001000000100",
"0000100000001000000000000000000000010100000000000000110000000001000000000110000000000010001000000100",
"0000100000001000000000000000000000010100000000000000110000000001000000000110000000000010001000000100",
"0000100000001000000000000000000000010100000000000000110000000001000000000110000000000010001000000100",
"0010101100000000110000000001010000011101000000100000110010001101100000010010100000000000001010100101",
"1101100010111110001011100010100100110100001110011010101101100011010011101110000110101011101001000100",
"1101100010001101001101100000101011101101001011011101101010110011011111101110000110111110001100111110",
"1101010010110010010101011101101111110110011000100110010000011000101000000101011110101110110001011111",
"0011001111111000001100100110100011000010101100110011000100010010010000100000101101101000101111001001",

"0000000100000100000000000010000000100000000000000000000000000000000000010000010000000000001000000000",
"0000000100000100000000000010000000100000000000000000000000000000000000010000010000000000001000000000",
"0000000100000100000000000010000000100000000000000000000000000000000000010000010000000000001000000000",
"0000000100000100000000000010000000100000000000000000000000000000000000010000010000000000001000000000",
"0000000100000100000000000010000000100000000000000000000000000000000000010000010000000000001000000000",
"0000000100000100000000000010000000100000000000000000000000000000000000010000010000000000001000000000",
"0001000101011010000100100000000000100101000000000000001001001001001010010000111000000100000001000000",
"0010001010100100011001001111101011000010111001011000110000110110110001001110000110100000001010011000",
"1100110010100101111001101010101101001000110111001000110100110110110000000101000001101001011010110100",
"1110010101000001011011010011111111101001111011110001011101110110000110101111110110011100110111111010",
"0110100011110101111000011010000001110000000001011111010110100100000111110111011110100110001000011111",

"0000010000010001000000100000000000000000000001000000000000010000000000000000000000000000000000000000",
"0000010000010001000000100000000000000000000001000000000000010000000000000000000000000000000000000000",
"0000010000010001000000100000000000000000000001000000000000010000000000000000000000000000000000000000",
"0000010000010001000000100000000000000000000001000000000000010000000000000000000000000000000000000000",
"0000010000010001000000100000000000000000000001000000000000010000000000000000000000000000000000000000",
"0000010000010001000000100000000000000000000001000000000000010000000000000000000000000000000000000000",
"1000010100101101110001100010000010000000010001000100000011110010001001000000000000001001110000011001",
"0000111001010010000000101001011100010111100000011011011000001001010100000111000000110100001110100110",
"0010010010011000101000001000000101100011101111010000001000110001110100001000101011110011001101100010",
"1111001100000110000011010010110011011010000111111011100100010100011110011110011110000000110100110110",
"1010111111110001000110010110101011101000011011011101100010011100010000101111110101001000101001110001",

"0000100000000000000010100110000000000000000000000000000000000000000000001010000000000000001101000000",
"0000100000000000000010100110000000000000000000000000000000000000000000001010000000000000001101000000",
"0000100000000000000010100110000000000000000000000000000000000000000000001010000000000000001101000000",
"0000100000000000000010100110000000000000000000000000000000000000000000001010000000000000001101000000",
"0000100000000000000010100110000000000000000000000000000000000000000000001010000000000000001101000000",
"0000100000000000000010100110000000000000000000000000000000000000000000001010000000000000001101000000",
"0001100100000001010110101100000100000011000000001000100000000010000100001010010000000001001101101000",
"1100000010111000000010010110001011001100000011110100010100001101010010111000001011110010001110010101",
"1010000011010110101001100010100010011000001000100110011001000100011001110101101100011110101010010111",
"0101011100100101110101110001010011100101101111000001001111111111100111010111110110001100111000100010",
"1010001100110010000000101000010101111100011011111001101000100000011110111011010011010001100010101101",

"0000000000000000000000000000000000000000000000000100100000100110010100010001001001001000010000001000",
"0000000000000000000000000000000000000000000000000100100000100110010100010001001001001000010000001000",
"0000000000000000000000000000000000000000000000000100100000100110010100010001001001001000010000001000",
"0000000000000000000000000000000000000000000000000100100000100110010100010001001001001000010000001000",
"0000000000000000000000000000000000000000000000000100100000100110010100010001001001001000010000001000",
"0000000000000000000000000000000000000000000000000100100000100110010100010001001001001000010000001000",
"0000010001000001000000010000101010000001000100000100100001100110110110011001011101001000011101001000",
"1001101110010010110111101111010001001100111011101110010110110001001101110100100011011110100000011100",
"1100000110011111001011000000010101100001001001010111001110111011011001010010111011001001000010001111",
"1111111110101010101110110100001010000000001110110100101110011000111011000100000001111000001101101110",
"1110001011101110010110100110100101011010100010110000011110111001000011001100101010110100011011000000",

"0000000000010000000000000000010000100000001000000000000000000000010000000000000000000000011000000000",
"0000000000010000000000000000010000100000001000000000000000000000010000000000000000000000011000000000",
"0000000000010000000000000000010000100000001000000000000000000000010000000000000000000000011000000000",
"0000000000010000000000000000010000100000001000000000000000000000010000000000000000000000011000000000",
"0000000000010000000000000000010000100000001000000000000000000000010000000000000000000000011000000000",
"0000000000010000000000000000010000100000001000000000000000000000010000000000000000000000011000000000",
"1000000000010001000000100100011000100110001000101101000000010001010000101001100000000001001010001000",
"0101000011001010101110011010110110011000010110010010100111000100010001010100011011101100110101100111",
"0011110001000111011011001001010011000001100100000010101100101110011110000000110001101010010100000000",
"0000101100111110110100100010010111110100010100110010010110101100110000010110011101111111001010111001",
"1110011111100010011100011111110001100000110011110100101000001000110111100001001111100001111011010110",

"0000000010000100000000000000000000000000010000000000001010000010000000000000000000000000100010000001",
"0000000010000100000000000000000000000000010000000000001010000010000000000000000000000000100010000001",
"0000000010000100000000000000000000000000010000000000001010000010000000000000000000000000100010000001",
"0000000010000100000000000000000000000000010000000000001010000010000000000000000000000000100010000001",
"0000000010000100000000000000000000000000010000000000001010000010000000000000000000000000100010000001",
"0000000010000100000000000000000000000000010000000000001010000010000000000000000000000000100010000001",
"0001001000011110000110000011001000000100000100100100000011000110010110000000000010011110100010001001",
"0010100110000100110001010100110110011011010010011000001000100011100000110011100001100001110101000100",
"0000110011110000001001011010010010110011010011001011011010111010101001101100110100110001011101100101",
"1110001110101101001100010001111101001001100100110111110111011001110101100000011101001111011110111001",
"1011001110100100110110101001101010000001011110111000001010111010000001101111010101100000110010001010",

"0000011000000000010000000000000000001100000000010000010100000000000001001000000001000000000110001000",
"0000011000000000010000000000000000001100000000010000010100000000000001001000000001000000000110001000",
"0000011000000000010000000000000000001100000000010000010100000000000001001000000001000000000110001000",
"0000011000000000010000000000000000001100000000010000010100000000000001001000000001000000000110001000",
"0000011000000000010000000000000000001100000000010000010100000000000001001000000001000000000110001000",
"0000011000000000010000000000000000001100000000010000010100000000000001001000000001000000000110001000",
"1000011000000010110111010000000100011000000010011000010111011000000001001000000000000100000110111001",
"0011100100011101001000101000100011100111101001000001101100100111001111011100010001010010000000001110",
"0010001011101101011010101001111011101101111101000101001000000100001001110101111101010010100001101010",
"0101111101100000101000100111100010110000011110011010110011001010110011000100001100100101101110011111",
"1110100001001000010100011101100001010101001001101101001001001111011101101110111111011010011001010011",

"0000001000000100000011000000000000001000000000100000000000000000000100010011000000000000000001000000",
"0000001000000100000011000000000000001000000000100000000000000000000100010011000000000000000001000000",
"0000001000000100000011000000000000001000000000100000000000000000000100010011000000000000000001000000",
"0000001000000100000011000000000000001000000000100000000000000000000100010011000000000000000001000000",
"0000001000000100000011000000000000001000000000100000000000000000000100010011000000000000000001000000",
"0000001000000100000011000000000000001000000000100000000000000000000100010011000000000000000001000000",
"1100101100000101000111001100100010101000001100101101000000010001101010010011000100000000000001000100",
"0011001010010010111010110001010000010011010010000000101001101000010101101111111011101111111011111011",
"0010111011110100001011100010001100000101110011010010101111000010010101011000101100110111111001001100",
"0110011110010011000011010000001101100001000001011100011011101110011010101010001001010000000100011011",
"0000001111101011111001000110111110101000000001001101001011100011110000111101101000101110110110001011"

);
end weight_mem_package;
package body weight_mem_package is
end weight_mem_package;
